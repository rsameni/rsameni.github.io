`ifndef _my_include_vh_
`define _my_include_vh_

`define W 700
`define DATA_LENGTH  16
`endif
