`timescale 1ns / 1ps
`include "macro.vh"
///////////////////////
module FIFO( in , out , clk ,reset);

input  [`DATA_LENGTH-1:0] in;
output [`DATA_LENGTH-1:0] out;
input  clk ,reset;
reg	[`DATA_LENGTH-1:0] fifo [0:`W-1];

assign  out =  fifo[`W-1] ;
always @(posedge clk)
begin
	if(reset)
	begin
		fifo[0] <= 0;
		fifo[1] <= 0;
		fifo[2] <= 0;
		fifo[3] <= 0;
		fifo[4] <= 0;
		fifo[5] <= 0;
		fifo[6] <= 0;
		fifo[7] <= 0;
		fifo[8] <= 0;
		fifo[9] <= 0;
		fifo[10] <= 0;
		fifo[11] <= 0;
		fifo[12] <= 0;
		fifo[13] <= 0;
		fifo[14] <= 0;
		fifo[15] <= 0;
		fifo[16] <= 0;
		fifo[17] <= 0;
		fifo[18] <= 0;
		fifo[19] <= 0;
		fifo[20] <= 0;
		fifo[21] <= 0;
		fifo[22] <= 0;
		fifo[23] <= 0;
		fifo[24] <= 0;
		fifo[25] <= 0;
		fifo[26] <= 0;
		fifo[27] <= 0;
		fifo[28] <= 0;
		fifo[29] <= 0;
		fifo[30] <= 0;
		fifo[31] <= 0;
		fifo[32] <= 0;
		fifo[33] <= 0;
		fifo[34] <= 0;
		fifo[35] <= 0;
		fifo[36] <= 0;
		fifo[37] <= 0;
		fifo[38] <= 0;
		fifo[39] <= 0;
		fifo[40] <= 0;
		fifo[41] <= 0;
		fifo[42] <= 0;
		fifo[43] <= 0;
		fifo[44] <= 0;
		fifo[45] <= 0;
		fifo[46] <= 0;
		fifo[47] <= 0;
		fifo[48] <= 0;
		fifo[49] <= 0;
		fifo[50] <= 0;
		fifo[51] <= 0;
		fifo[52] <= 0;
		fifo[53] <= 0;
		fifo[54] <= 0;
		fifo[55] <= 0;
		fifo[56] <= 0;
		fifo[57] <= 0;
		fifo[58] <= 0;
		fifo[59] <= 0;
		fifo[60] <= 0;
		fifo[61] <= 0;
		fifo[62] <= 0;
		fifo[63] <= 0;
		fifo[64] <= 0;
		fifo[65] <= 0;
		fifo[66] <= 0;
		fifo[67] <= 0;
		fifo[68] <= 0;
		fifo[69] <= 0;
		fifo[70] <= 0;
		fifo[71] <= 0;
		fifo[72] <= 0;
		fifo[73] <= 0;
		fifo[74] <= 0;
		fifo[75] <= 0;
		fifo[76] <= 0;
		fifo[77] <= 0;
		fifo[78] <= 0;
		fifo[79] <= 0;
		fifo[80] <= 0;
		fifo[81] <= 0;
		fifo[82] <= 0;
		fifo[83] <= 0;
		fifo[84] <= 0;
		fifo[85] <= 0;
		fifo[86] <= 0;
		fifo[87] <= 0;
		fifo[88] <= 0;
		fifo[89] <= 0;
		fifo[90] <= 0;
		fifo[91] <= 0;
		fifo[92] <= 0;
		fifo[93] <= 0;
		fifo[94] <= 0;
		fifo[95] <= 0;
		fifo[96] <= 0;
		fifo[97] <= 0;
		fifo[98] <= 0;
		fifo[99] <= 0;
		fifo[100] <= 0;
		fifo[101] <= 0;
		fifo[102] <= 0;
		fifo[103] <= 0;
		fifo[104] <= 0;
		fifo[105] <= 0;
		fifo[106] <= 0;
		fifo[107] <= 0;
		fifo[108] <= 0;
		fifo[109] <= 0;
		fifo[110] <= 0;
		fifo[111] <= 0;
		fifo[112] <= 0;
		fifo[113] <= 0;
		fifo[114] <= 0;
		fifo[115] <= 0;
		fifo[116] <= 0;
		fifo[117] <= 0;
		fifo[118] <= 0;
		fifo[119] <= 0;
		fifo[120] <= 0;
		fifo[121] <= 0;
		fifo[122] <= 0;
		fifo[123] <= 0;
		fifo[124] <= 0;
		fifo[125] <= 0;
		fifo[126] <= 0;
		fifo[127] <= 0;
		fifo[128] <= 0;
		fifo[129] <= 0;
		fifo[130] <= 0;
		fifo[131] <= 0;
		fifo[132] <= 0;
		fifo[133] <= 0;
		fifo[134] <= 0;
		fifo[135] <= 0;
		fifo[136] <= 0;
		fifo[137] <= 0;
		fifo[138] <= 0;
		fifo[139] <= 0;
		fifo[140] <= 0;
		fifo[141] <= 0;
		fifo[142] <= 0;
		fifo[143] <= 0;
		fifo[144] <= 0;
		fifo[145] <= 0;
		fifo[146] <= 0;
		fifo[147] <= 0;
		fifo[148] <= 0;
		fifo[149] <= 0;
		fifo[150] <= 0;
		fifo[151] <= 0;
		fifo[152] <= 0;
		fifo[153] <= 0;
		fifo[154] <= 0;
		fifo[155] <= 0;
		fifo[156] <= 0;
		fifo[157] <= 0;
		fifo[158] <= 0;
		fifo[159] <= 0;
		fifo[160] <= 0;
		fifo[161] <= 0;
		fifo[162] <= 0;
		fifo[163] <= 0;
		fifo[164] <= 0;
		fifo[165] <= 0;
		fifo[166] <= 0;
		fifo[167] <= 0;
		fifo[168] <= 0;
		fifo[169] <= 0;
		fifo[170] <= 0;
		fifo[171] <= 0;
		fifo[172] <= 0;
		fifo[173] <= 0;
		fifo[174] <= 0;
		fifo[175] <= 0;
		fifo[176] <= 0;
		fifo[177] <= 0;
		fifo[178] <= 0;
		fifo[179] <= 0;
		fifo[180] <= 0;
		fifo[181] <= 0;
		fifo[182] <= 0;
		fifo[183] <= 0;
		fifo[184] <= 0;
		fifo[185] <= 0;
		fifo[186] <= 0;
		fifo[187] <= 0;
		fifo[188] <= 0;
		fifo[189] <= 0;
		fifo[190] <= 0;
		fifo[191] <= 0;
		fifo[192] <= 0;
		fifo[193] <= 0;
		fifo[194] <= 0;
		fifo[195] <= 0;
		fifo[196] <= 0;
		fifo[197] <= 0;
		fifo[198] <= 0;
		fifo[199] <= 0;
		fifo[200] <= 0;
		fifo[201] <= 0;
		fifo[202] <= 0;
		fifo[203] <= 0;
		fifo[204] <= 0;
		fifo[205] <= 0;
		fifo[206] <= 0;
		fifo[207] <= 0;
		fifo[208] <= 0;
		fifo[209] <= 0;
		fifo[210] <= 0;
		fifo[211] <= 0;
		fifo[212] <= 0;
		fifo[213] <= 0;
		fifo[214] <= 0;
		fifo[215] <= 0;
		fifo[216] <= 0;
		fifo[217] <= 0;
		fifo[218] <= 0;
		fifo[219] <= 0;
		fifo[220] <= 0;
		fifo[221] <= 0;
		fifo[222] <= 0;
		fifo[223] <= 0;
		fifo[224] <= 0;
		fifo[225] <= 0;
		fifo[226] <= 0;
		fifo[227] <= 0;
		fifo[228] <= 0;
		fifo[229] <= 0;
		fifo[230] <= 0;
		fifo[231] <= 0;
		fifo[232] <= 0;
		fifo[233] <= 0;
		fifo[234] <= 0;
		fifo[235] <= 0;
		fifo[236] <= 0;
		fifo[237] <= 0;
		fifo[238] <= 0;
		fifo[239] <= 0;
		fifo[240] <= 0;
		fifo[241] <= 0;
		fifo[242] <= 0;
		fifo[243] <= 0;
		fifo[244] <= 0;
		fifo[245] <= 0;
		fifo[246] <= 0;
		fifo[247] <= 0;
		fifo[248] <= 0;
		fifo[249] <= 0;
		fifo[250] <= 0;
		fifo[251] <= 0;
		fifo[252] <= 0;
		fifo[253] <= 0;
		fifo[254] <= 0;
		fifo[255] <= 0;
		fifo[256] <= 0;
		fifo[257] <= 0;
		fifo[258] <= 0;
		fifo[259] <= 0;
		fifo[260] <= 0;
		fifo[261] <= 0;
		fifo[262] <= 0;
		fifo[263] <= 0;
		fifo[264] <= 0;
		fifo[265] <= 0;
		fifo[266] <= 0;
		fifo[267] <= 0;
		fifo[268] <= 0;
		fifo[269] <= 0;
		fifo[270] <= 0;
		fifo[271] <= 0;
		fifo[272] <= 0;
		fifo[273] <= 0;
		fifo[274] <= 0;
		fifo[275] <= 0;
		fifo[276] <= 0;
		fifo[277] <= 0;
		fifo[278] <= 0;
		fifo[279] <= 0;
		fifo[280] <= 0;
		fifo[281] <= 0;
		fifo[282] <= 0;
		fifo[283] <= 0;
		fifo[284] <= 0;
		fifo[285] <= 0;
		fifo[286] <= 0;
		fifo[287] <= 0;
		fifo[288] <= 0;
		fifo[289] <= 0;
		fifo[290] <= 0;
		fifo[291] <= 0;
		fifo[292] <= 0;
		fifo[293] <= 0;
		fifo[294] <= 0;
		fifo[295] <= 0;
		fifo[296] <= 0;
		fifo[297] <= 0;
		fifo[298] <= 0;
		fifo[299] <= 0;
	end
	else
	begin
			fifo[0] <= in ;
			fifo[1] <= fifo[0];
			fifo[2] <= fifo[1];
			fifo[3] <= fifo[2];
			fifo[4] <= fifo[3];
			fifo[5] <= fifo[4];
			fifo[6] <= fifo[5];
			fifo[7] <= fifo[6];
			fifo[8] <= fifo[7];
			fifo[9] <= fifo[8];
			fifo[10] <= fifo[9];
			fifo[11] <= fifo[10];
			fifo[12] <= fifo[11];
			fifo[13] <= fifo[12];
			fifo[14] <= fifo[13];
			fifo[15] <= fifo[14];
			fifo[16] <= fifo[15];
			fifo[17] <= fifo[16];
			fifo[18] <= fifo[17];
			fifo[19] <= fifo[18];
			fifo[20] <= fifo[19];
			fifo[21] <= fifo[20];
			fifo[22] <= fifo[21];
			fifo[23] <= fifo[22];
			fifo[24] <= fifo[23];
			fifo[25] <= fifo[24];
			fifo[26] <= fifo[25];
			fifo[27] <= fifo[26];
			fifo[28] <= fifo[27];
			fifo[29] <= fifo[28];
			fifo[30] <= fifo[29];
			fifo[31] <= fifo[30];
			fifo[32] <= fifo[31];
			fifo[33] <= fifo[32];
			fifo[34] <= fifo[33];
			fifo[35] <= fifo[34];
			fifo[36] <= fifo[35];
			fifo[37] <= fifo[36];
			fifo[38] <= fifo[37];
			fifo[39] <= fifo[38];
			fifo[40] <= fifo[39];
			fifo[41] <= fifo[40];
			fifo[42] <= fifo[41];
			fifo[43] <= fifo[42];
			fifo[44] <= fifo[43];
			fifo[45] <= fifo[44];
			fifo[46] <= fifo[45];
			fifo[47] <= fifo[46];
			fifo[48] <= fifo[47];
			fifo[49] <= fifo[48];
			fifo[50] <= fifo[49];
			fifo[51] <= fifo[50];
			fifo[52] <= fifo[51];
			fifo[53] <= fifo[52];
			fifo[54] <= fifo[53];
			fifo[55] <= fifo[54];
			fifo[56] <= fifo[55];
			fifo[57] <= fifo[56];
			fifo[58] <= fifo[57];
			fifo[59] <= fifo[58];
			fifo[60] <= fifo[59];
			fifo[61] <= fifo[60];
			fifo[62] <= fifo[61];
			fifo[63] <= fifo[62];
			fifo[64] <= fifo[63];
			fifo[65] <= fifo[64];
			fifo[66] <= fifo[65];
			fifo[67] <= fifo[66];
			fifo[68] <= fifo[67];
			fifo[69] <= fifo[68];
			fifo[70] <= fifo[69];
			fifo[71] <= fifo[70];
			fifo[72] <= fifo[71];
			fifo[73] <= fifo[72];
			fifo[74] <= fifo[73];
			fifo[75] <= fifo[74];
			fifo[76] <= fifo[75];
			fifo[77] <= fifo[76];
			fifo[78] <= fifo[77];
			fifo[79] <= fifo[78];
			fifo[80] <= fifo[79];
			fifo[81] <= fifo[80];
			fifo[82] <= fifo[81];
			fifo[83] <= fifo[82];
			fifo[84] <= fifo[83];
			fifo[85] <= fifo[84];
			fifo[86] <= fifo[85];
			fifo[87] <= fifo[86];
			fifo[88] <= fifo[87];
			fifo[89] <= fifo[88];
			fifo[90] <= fifo[89];
			fifo[91] <= fifo[90];
			fifo[92] <= fifo[91];
			fifo[93] <= fifo[92];
			fifo[94] <= fifo[93];
			fifo[95] <= fifo[94];
			fifo[96] <= fifo[95];
			fifo[97] <= fifo[96];
			fifo[98] <= fifo[97];
			fifo[99] <= fifo[98];
			fifo[100] <= fifo[99];
			fifo[101] <= fifo[100];
			fifo[102] <= fifo[101];
			fifo[103] <= fifo[102];
			fifo[104] <= fifo[103];
			fifo[105] <= fifo[104];
			fifo[106] <= fifo[105];
			fifo[107] <= fifo[106];
			fifo[108] <= fifo[107];
			fifo[109] <= fifo[108];
			fifo[110] <= fifo[109];
			fifo[111] <= fifo[110];
			fifo[112] <= fifo[111];
			fifo[113] <= fifo[112];
			fifo[114] <= fifo[113];
			fifo[115] <= fifo[114];
			fifo[116] <= fifo[115];
			fifo[117] <= fifo[116];
			fifo[118] <= fifo[117];
			fifo[119] <= fifo[118];
			fifo[120] <= fifo[119];
			fifo[121] <= fifo[120];
			fifo[122] <= fifo[121];
			fifo[123] <= fifo[122];
			fifo[124] <= fifo[123];
			fifo[125] <= fifo[124];
			fifo[126] <= fifo[125];
			fifo[127] <= fifo[126];
			fifo[128] <= fifo[127];
			fifo[129] <= fifo[128];
			fifo[130] <= fifo[129];
			fifo[131] <= fifo[130];
			fifo[132] <= fifo[131];
			fifo[133] <= fifo[132];
			fifo[134] <= fifo[133];
			fifo[135] <= fifo[134];
			fifo[136] <= fifo[135];
			fifo[137] <= fifo[136];
			fifo[138] <= fifo[137];
			fifo[139] <= fifo[138];
			fifo[140] <= fifo[139];
			fifo[141] <= fifo[140];
			fifo[142] <= fifo[141];
			fifo[143] <= fifo[142];
			fifo[144] <= fifo[143];
			fifo[145] <= fifo[144];
			fifo[146] <= fifo[145];
			fifo[147] <= fifo[146];
			fifo[148] <= fifo[147];
			fifo[149] <= fifo[148];
			fifo[150] <= fifo[149];
			fifo[151] <= fifo[150];
			fifo[152] <= fifo[151];
			fifo[153] <= fifo[152];
			fifo[154] <= fifo[153];
			fifo[155] <= fifo[154];
			fifo[156] <= fifo[155];
			fifo[157] <= fifo[156];
			fifo[158] <= fifo[157];
			fifo[159] <= fifo[158];
			fifo[160] <= fifo[159];
			fifo[161] <= fifo[160];
			fifo[162] <= fifo[161];
			fifo[163] <= fifo[162];
			fifo[164] <= fifo[163];
			fifo[165] <= fifo[164];
			fifo[166] <= fifo[165];
			fifo[167] <= fifo[166];
			fifo[168] <= fifo[167];
			fifo[169] <= fifo[168];
			fifo[170] <= fifo[169];
			fifo[171] <= fifo[170];
			fifo[172] <= fifo[171];
			fifo[173] <= fifo[172];
			fifo[174] <= fifo[173];
			fifo[175] <= fifo[174];
			fifo[176] <= fifo[175];
			fifo[177] <= fifo[176];
			fifo[178] <= fifo[177];
			fifo[179] <= fifo[178];
			fifo[180] <= fifo[179];
			fifo[181] <= fifo[180];
			fifo[182] <= fifo[181];
			fifo[183] <= fifo[182];
			fifo[184] <= fifo[183];
			fifo[185] <= fifo[184];
			fifo[186] <= fifo[185];
			fifo[187] <= fifo[186];
			fifo[188] <= fifo[187];
			fifo[189] <= fifo[188];
			fifo[190] <= fifo[189];
			fifo[191] <= fifo[190];
			fifo[192] <= fifo[191];
			fifo[193] <= fifo[192];
			fifo[194] <= fifo[193];
			fifo[195] <= fifo[194];
			fifo[196] <= fifo[195];
			fifo[197] <= fifo[196];
			fifo[198] <= fifo[197];
			fifo[199] <= fifo[198];
			fifo[200] <= fifo[199];
			fifo[201] <= fifo[200];
			fifo[202] <= fifo[201];
			fifo[203] <= fifo[202];
			fifo[204] <= fifo[203];
			fifo[205] <= fifo[204];
			fifo[206] <= fifo[205];
			fifo[207] <= fifo[206];
			fifo[208] <= fifo[207];
			fifo[209] <= fifo[208];
			fifo[210] <= fifo[209];
			fifo[211] <= fifo[210];
			fifo[212] <= fifo[211];
			fifo[213] <= fifo[212];
			fifo[214] <= fifo[213];
			fifo[215] <= fifo[214];
			fifo[216] <= fifo[215];
			fifo[217] <= fifo[216];
			fifo[218] <= fifo[217];
			fifo[219] <= fifo[218];
			fifo[220] <= fifo[219];
			fifo[221] <= fifo[220];
			fifo[222] <= fifo[221];
			fifo[223] <= fifo[222];
			fifo[224] <= fifo[223];
			fifo[225] <= fifo[224];
			fifo[226] <= fifo[225];
			fifo[227] <= fifo[226];
			fifo[228] <= fifo[227];
			fifo[229] <= fifo[228];
			fifo[230] <= fifo[229];
			fifo[231] <= fifo[230];
			fifo[232] <= fifo[231];
			fifo[233] <= fifo[232];
			fifo[234] <= fifo[233];
			fifo[235] <= fifo[234];
			fifo[236] <= fifo[235];
			fifo[237] <= fifo[236];
			fifo[238] <= fifo[237];
			fifo[239] <= fifo[238];
			fifo[240] <= fifo[239];
			fifo[241] <= fifo[240];
			fifo[242] <= fifo[241];
			fifo[243] <= fifo[242];
			fifo[244] <= fifo[243];
			fifo[245] <= fifo[244];
			fifo[246] <= fifo[245];
			fifo[247] <= fifo[246];
			fifo[248] <= fifo[247];
			fifo[249] <= fifo[248];
			fifo[250] <= fifo[249];
			fifo[251] <= fifo[250];
			fifo[252] <= fifo[251];
			fifo[253] <= fifo[252];
			fifo[254] <= fifo[253];
			fifo[255] <= fifo[254];
			fifo[256] <= fifo[255];
			fifo[257] <= fifo[256];
			fifo[258] <= fifo[257];
			fifo[259] <= fifo[258];
			fifo[260] <= fifo[259];
			fifo[261] <= fifo[260];
			fifo[262] <= fifo[261];
			fifo[263] <= fifo[262];
			fifo[264] <= fifo[263];
			fifo[265] <= fifo[264];
			fifo[266] <= fifo[265];
			fifo[267] <= fifo[266];
			fifo[268] <= fifo[267];
			fifo[269] <= fifo[268];
			fifo[270] <= fifo[269];
			fifo[271] <= fifo[270];
			fifo[272] <= fifo[271];
			fifo[273] <= fifo[272];
			fifo[274] <= fifo[273];
			fifo[275] <= fifo[274];
			fifo[276] <= fifo[275];
			fifo[277] <= fifo[276];
			fifo[278] <= fifo[277];
			fifo[279] <= fifo[278];
			fifo[280] <= fifo[279];
			fifo[281] <= fifo[280];
			fifo[282] <= fifo[281];
			fifo[283] <= fifo[282];
			fifo[284] <= fifo[283];
			fifo[285] <= fifo[284];
			fifo[286] <= fifo[285];
			fifo[287] <= fifo[286];
			fifo[288] <= fifo[287];
			fifo[289] <= fifo[288];
			fifo[290] <= fifo[289];
			fifo[291] <= fifo[290];
			fifo[292] <= fifo[291];
			fifo[293] <= fifo[292];
			fifo[294] <= fifo[293];
			fifo[295] <= fifo[294];
			fifo[296] <= fifo[295];
			fifo[297] <= fifo[296];
			fifo[298] <= fifo[297];
			fifo[299] <= fifo[298];
	end
end

endmodule