`ifndef _my_include_vh_
`define _my_include_vh_

`define W_MAX 201
`define LOG_WMAX 8
`define DATA_LENGTH  16
`define HIGH_Z  16'bz
`endif
