`timescale 1ns / 1ps
`include "macro.vh"
///////////////////////
module top ( clk ,reset ,X ,median );

output [`DATA_LENGTH-1:0] median ;
input [`DATA_LENGTH-1:0] X ;
input clk ,reset ;

wire 	[`DATA_LENGTH-1:0] R_old, R1 ,R2 ,R3 ,R4 ,R5 ,R6 ,R7 ,R8 ,R9 ,R10 ,R11 ,R12 ,R13 ,R14 ,R15 ,R16 ,R17 ,R18 ,R19 ,R20 ,R21 ,R22 ,R23 ,R24 ,R25 ,R26 ,R27 ,R28 ,R29 ,R30 ,R31 ,R32 ,R33 ,R34 ,R35 ,R36 ,R37 ,R38 ,R39 ,R40 ,R41 ,R42 ,R43 ,R44 ,R45 ,R46 ,R47 ,R48 ,R49 ,R50 ,R51 ,R52 ,R53 ,R54 ,R55 ,R56 ,R57 ,R58 ,R59 ,R60 ,R61 ,R62 ,R63 ,R64 ,R65 ,R66 ,R67 ,R68 ,R69 ,R70 ,R71 ,R72 ,R73 ,R74 ,R75 ,R76 ,R77 ,R78 ,R79 ,R80 ,R81 ,R82 ,R83 ,R84 ,R85 ,R86 ,R87 ,R88 ,R89 ,R90 ,R91 ,R92 ,R93 ,R94 ,R95 ,R96 ,R97 ,R98 ,R99 ,R100 ,R101 ,R102 ,R103 ,R104 ,R105 ,R106 ,R107 ,R108 ,R109 ,R110 ,R111 ,R112 ,R113 ,R114 ,R115 ,R116 ,R117 ,R118 ,R119 ,R120 ,R121 ,R122 ,R123 ,R124 ,R125 ,R126 ,R127 ,R128 ,R129 ,R130 ,R131 ,R132 ,R133 ,R134 ,R135 ,R136 ,R137 ,R138 ,R139 ,R140 ,R141 ,R142 ,R143 ,R144 ,R145 ,R146 ,R147 ,R148 ,R149 ,R150 ,R151 ,R152 ,R153 ,R154 ,R155 ,R156 ,R157 ,R158 ,R159 ,R160 ,R161 ,R162 ,R163 ,R164 ,R165 ,R166 ,R167 ,R168 ,R169 ,R170 ,R171 ,R172 ,R173 ,R174 ,R175 ,R176 ,R177 ,R178 ,R179 ,R180 ,R181 ,R182 ,R183 ,R184 ,R185 ,R186 ,R187 ,R188 ,R189 ,R190 ,R191 ,R192 ,R193 ,R194 ,R195 ,R196 ,R197 ,R198 ,R199 ,R200 ,R201 ,R202 ,R203 ,R204 ,R205 ,R206 ,R207 ,R208 ,R209 ,R210 ,R211 ,R212 ,R213 ,R214 ,R215 ,R216 ,R217 ,R218 ,R219 ,R220 ,R221 ,R222 ,R223 ,R224 ,R225 ,R226 ,R227 ,R228 ,R229 ,R230 ,R231 ,R232 ,R233 ,R234 ,R235 ,R236 ,R237 ,R238 ,R239 ,R240 ,R241 ,R242 ,R243 ,R244 ,R245 ,R246 ,R247 ,R248 ,R249 ,R250 ,R251 ,R252 ,R253 ,R254 ,R255 ,R256 ,R257 ,R258 ,R259 ,R260 ,R261 ,R262 ,R263 ,R264 ,R265 ,R266 ,R267 ,R268 ,R269 ,R270 ,R271 ,R272 ,R273 ,R274 ,R275 ,R276 ,R277 ,R278 ,R279 ,R280 ,R281 ,R282 ,R283 ,R284 ,R285 ,R286 ,R287 ,R288 ,R289 ,R290 ,R291 ,R292 ,R293 ,R294 ,R295 ,R296 ,R297 ,R298 ,R299 ,R300;
wire 	T1 ,T2 ,T3 ,T4 ,T5 ,T6 ,T7 ,T8 ,T9 ,T10 ,T11 ,T12 ,T13 ,T14 ,T15 ,T16 ,T17 ,T18 ,T19 ,T20 ,T21 ,T22 ,T23 ,T24 ,T25 ,T26 ,T27 ,T28 ,T29 ,T30 ,T31 ,T32 ,T33 ,T34 ,T35 ,T36 ,T37 ,T38 ,T39 ,T40 ,T41 ,T42 ,T43 ,T44 ,T45 ,T46 ,T47 ,T48 ,T49 ,T50 ,T51 ,T52 ,T53 ,T54 ,T55 ,T56 ,T57 ,T58 ,T59 ,T60 ,T61 ,T62 ,T63 ,T64 ,T65 ,T66 ,T67 ,T68 ,T69 ,T70 ,T71 ,T72 ,T73 ,T74 ,T75 ,T76 ,T77 ,T78 ,T79 ,T80 ,T81 ,T82 ,T83 ,T84 ,T85 ,T86 ,T87 ,T88 ,T89 ,T90 ,T91 ,T92 ,T93 ,T94 ,T95 ,T96 ,T97 ,T98 ,T99 ,T100 ,T101 ,T102 ,T103 ,T104 ,T105 ,T106 ,T107 ,T108 ,T109 ,T110 ,T111 ,T112 ,T113 ,T114 ,T115 ,T116 ,T117 ,T118 ,T119 ,T120 ,T121 ,T122 ,T123 ,T124 ,T125 ,T126 ,T127 ,T128 ,T129 ,T130 ,T131 ,T132 ,T133 ,T134 ,T135 ,T136 ,T137 ,T138 ,T139 ,T140 ,T141 ,T142 ,T143 ,T144 ,T145 ,T146 ,T147 ,T148 ,T149 ,T150 ,T151 ,T152 ,T153 ,T154 ,T155 ,T156 ,T157 ,T158 ,T159 ,T160 ,T161 ,T162 ,T163 ,T164 ,T165 ,T166 ,T167 ,T168 ,T169 ,T170 ,T171 ,T172 ,T173 ,T174 ,T175 ,T176 ,T177 ,T178 ,T179 ,T180 ,T181 ,T182 ,T183 ,T184 ,T185 ,T186 ,T187 ,T188 ,T189 ,T190 ,T191 ,T192 ,T193 ,T194 ,T195 ,T196 ,T197 ,T198 ,T199 ,T200 ,T201 ,T202 ,T203 ,T204 ,T205 ,T206 ,T207 ,T208 ,T209 ,T210 ,T211 ,T212 ,T213 ,T214 ,T215 ,T216 ,T217 ,T218 ,T219 ,T220 ,T221 ,T222 ,T223 ,T224 ,T225 ,T226 ,T227 ,T228 ,T229 ,T230 ,T231 ,T232 ,T233 ,T234 ,T235 ,T236 ,T237 ,T238 ,T239 ,T240 ,T241 ,T242 ,T243 ,T244 ,T245 ,T246 ,T247 ,T248 ,T249 ,T250 ,T251 ,T252 ,T253 ,T254 ,T255 ,T256 ,T257 ,T258 ,T259 ,T260 ,T261 ,T262 ,T263 ,T264 ,T265 ,T266 ,T267 ,T268 ,T269 ,T270 ,T271 ,T272 ,T273 ,T274 ,T275 ,T276 ,T277 ,T278 ,T279 ,T280 ,T281 ,T282 ,T283 ,T284 ,T285 ,T286 ,T287 ,T288 ,T289 ,T290 ,T291 ,T292 ,T293 ,T294 ,T295 ,T296 ,T297 ,T298 ,T299 ,T300;
wire 	 Z1 ,Z2 ,Z3 ,Z4 ,Z5 ,Z6 ,Z7 ,Z8 ,Z9 ,Z10 ,Z11 ,Z12 ,Z13 ,Z14 ,Z15 ,Z16 ,Z17 ,Z18 ,Z19 ,Z20 ,Z21 ,Z22 ,Z23 ,Z24 ,Z25 ,Z26 ,Z27 ,Z28 ,Z29 ,Z30 ,Z31 ,Z32 ,Z33 ,Z34 ,Z35 ,Z36 ,Z37 ,Z38 ,Z39 ,Z40 ,Z41 ,Z42 ,Z43 ,Z44 ,Z45 ,Z46 ,Z47 ,Z48 ,Z49 ,Z50 ,Z51 ,Z52 ,Z53 ,Z54 ,Z55 ,Z56 ,Z57 ,Z58 ,Z59 ,Z60 ,Z61 ,Z62 ,Z63 ,Z64 ,Z65 ,Z66 ,Z67 ,Z68 ,Z69 ,Z70 ,Z71 ,Z72 ,Z73 ,Z74 ,Z75 ,Z76 ,Z77 ,Z78 ,Z79 ,Z80 ,Z81 ,Z82 ,Z83 ,Z84 ,Z85 ,Z86 ,Z87 ,Z88 ,Z89 ,Z90 ,Z91 ,Z92 ,Z93 ,Z94 ,Z95 ,Z96 ,Z97 ,Z98 ,Z99 ,Z100 ,Z101 ,Z102 ,Z103 ,Z104 ,Z105 ,Z106 ,Z107 ,Z108 ,Z109 ,Z110 ,Z111 ,Z112 ,Z113 ,Z114 ,Z115 ,Z116 ,Z117 ,Z118 ,Z119 ,Z120 ,Z121 ,Z122 ,Z123 ,Z124 ,Z125 ,Z126 ,Z127 ,Z128 ,Z129 ,Z130 ,Z131 ,Z132 ,Z133 ,Z134 ,Z135 ,Z136 ,Z137 ,Z138 ,Z139 ,Z140 ,Z141 ,Z142 ,Z143 ,Z144 ,Z145 ,Z146 ,Z147 ,Z148 ,Z149 ,Z150 ,Z151 ,Z152 ,Z153 ,Z154 ,Z155 ,Z156 ,Z157 ,Z158 ,Z159 ,Z160 ,Z161 ,Z162 ,Z163 ,Z164 ,Z165 ,Z166 ,Z167 ,Z168 ,Z169 ,Z170 ,Z171 ,Z172 ,Z173 ,Z174 ,Z175 ,Z176 ,Z177 ,Z178 ,Z179 ,Z180 ,Z181 ,Z182 ,Z183 ,Z184 ,Z185 ,Z186 ,Z187 ,Z188 ,Z189 ,Z190 ,Z191 ,Z192 ,Z193 ,Z194 ,Z195 ,Z196 ,Z197 ,Z198 ,Z199 ,Z200 ,Z201 ,Z202 ,Z203 ,Z204 ,Z205 ,Z206 ,Z207 ,Z208 ,Z209 ,Z210 ,Z211 ,Z212 ,Z213 ,Z214 ,Z215 ,Z216 ,Z217 ,Z218 ,Z219 ,Z220 ,Z221 ,Z222 ,Z223 ,Z224 ,Z225 ,Z226 ,Z227 ,Z228 ,Z229 ,Z230 ,Z231 ,Z232 ,Z233 ,Z234 ,Z235 ,Z236 ,Z237 ,Z238 ,Z239 ,Z240 ,Z241 ,Z242 ,Z243 ,Z244 ,Z245 ,Z246 ,Z247 ,Z248 ,Z249 ,Z250 ,Z251 ,Z252 ,Z253 ,Z254 ,Z255 ,Z256 ,Z257 ,Z258 ,Z259 ,Z260 ,Z261 ,Z262 ,Z263 ,Z264 ,Z265 ,Z266 ,Z267 ,Z268 ,Z269 ,Z270 ,Z271 ,Z272 ,Z273 ,Z274 ,Z275 ,Z276 ,Z277 ,Z278 ,Z279 ,Z280 ,Z281 ,Z282 ,Z283 ,Z284 ,Z285 ,Z286 ,Z287 ,Z288 ,Z289 ,Z290 ,Z291 ,Z292 ,Z293 ,Z294 ,Z295 ,Z296 ,Z297 ,Z298 ,Z299;
 assign median = (R150 + R151)>>1;

FIFO myfifo(.in(X), .out(R_old), .clk(clk), .reset(reset));
medianCell_leftMst  m1(.X(X) , .clk(clk), .reset(reset) , .R_R(R2), .T_R(T2), .R_old(R_old), .Z(Z1), .R(R1), .T(T1));
medianFilterCell  m2(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z1), .R_L(R1),.R_R(R3) ,.T_L(T1), .T_R(T3), .R_old(R_old), .Z(Z2), .R(R2), .T(T2));
medianFilterCell  m3(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z2), .R_L(R2),.R_R(R4) ,.T_L(T2), .T_R(T4), .R_old(R_old), .Z(Z3), .R(R3), .T(T3));
medianFilterCell  m4(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z3), .R_L(R3),.R_R(R5) ,.T_L(T3), .T_R(T5), .R_old(R_old), .Z(Z4), .R(R4), .T(T4));
medianFilterCell  m5(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z4), .R_L(R4),.R_R(R6) ,.T_L(T4), .T_R(T6), .R_old(R_old), .Z(Z5), .R(R5), .T(T5));
medianFilterCell  m6(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z5), .R_L(R5),.R_R(R7) ,.T_L(T5), .T_R(T7), .R_old(R_old), .Z(Z6), .R(R6), .T(T6));
medianFilterCell  m7(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z6), .R_L(R6),.R_R(R8) ,.T_L(T6), .T_R(T8), .R_old(R_old), .Z(Z7), .R(R7), .T(T7));
medianFilterCell  m8(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z7), .R_L(R7),.R_R(R9) ,.T_L(T7), .T_R(T9), .R_old(R_old), .Z(Z8), .R(R8), .T(T8));
medianFilterCell  m9(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z8), .R_L(R8),.R_R(R10) ,.T_L(T8), .T_R(T10), .R_old(R_old), .Z(Z9), .R(R9), .T(T9));
medianFilterCell  m10(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z9), .R_L(R9),.R_R(R11) ,.T_L(T9), .T_R(T11), .R_old(R_old), .Z(Z10), .R(R10), .T(T10));
medianFilterCell  m11(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z10), .R_L(R10),.R_R(R12) ,.T_L(T10), .T_R(T12), .R_old(R_old), .Z(Z11), .R(R11), .T(T11));
medianFilterCell  m12(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z11), .R_L(R11),.R_R(R13) ,.T_L(T11), .T_R(T13), .R_old(R_old), .Z(Z12), .R(R12), .T(T12));
medianFilterCell  m13(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z12), .R_L(R12),.R_R(R14) ,.T_L(T12), .T_R(T14), .R_old(R_old), .Z(Z13), .R(R13), .T(T13));
medianFilterCell  m14(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z13), .R_L(R13),.R_R(R15) ,.T_L(T13), .T_R(T15), .R_old(R_old), .Z(Z14), .R(R14), .T(T14));
medianFilterCell  m15(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z14), .R_L(R14),.R_R(R16) ,.T_L(T14), .T_R(T16), .R_old(R_old), .Z(Z15), .R(R15), .T(T15));
medianFilterCell  m16(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z15), .R_L(R15),.R_R(R17) ,.T_L(T15), .T_R(T17), .R_old(R_old), .Z(Z16), .R(R16), .T(T16));
medianFilterCell  m17(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z16), .R_L(R16),.R_R(R18) ,.T_L(T16), .T_R(T18), .R_old(R_old), .Z(Z17), .R(R17), .T(T17));
medianFilterCell  m18(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z17), .R_L(R17),.R_R(R19) ,.T_L(T17), .T_R(T19), .R_old(R_old), .Z(Z18), .R(R18), .T(T18));
medianFilterCell  m19(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z18), .R_L(R18),.R_R(R20) ,.T_L(T18), .T_R(T20), .R_old(R_old), .Z(Z19), .R(R19), .T(T19));
medianFilterCell  m20(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z19), .R_L(R19),.R_R(R21) ,.T_L(T19), .T_R(T21), .R_old(R_old), .Z(Z20), .R(R20), .T(T20));
medianFilterCell  m21(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z20), .R_L(R20),.R_R(R22) ,.T_L(T20), .T_R(T22), .R_old(R_old), .Z(Z21), .R(R21), .T(T21));
medianFilterCell  m22(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z21), .R_L(R21),.R_R(R23) ,.T_L(T21), .T_R(T23), .R_old(R_old), .Z(Z22), .R(R22), .T(T22));
medianFilterCell  m23(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z22), .R_L(R22),.R_R(R24) ,.T_L(T22), .T_R(T24), .R_old(R_old), .Z(Z23), .R(R23), .T(T23));
medianFilterCell  m24(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z23), .R_L(R23),.R_R(R25) ,.T_L(T23), .T_R(T25), .R_old(R_old), .Z(Z24), .R(R24), .T(T24));
medianFilterCell  m25(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z24), .R_L(R24),.R_R(R26) ,.T_L(T24), .T_R(T26), .R_old(R_old), .Z(Z25), .R(R25), .T(T25));
medianFilterCell  m26(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z25), .R_L(R25),.R_R(R27) ,.T_L(T25), .T_R(T27), .R_old(R_old), .Z(Z26), .R(R26), .T(T26));
medianFilterCell  m27(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z26), .R_L(R26),.R_R(R28) ,.T_L(T26), .T_R(T28), .R_old(R_old), .Z(Z27), .R(R27), .T(T27));
medianFilterCell  m28(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z27), .R_L(R27),.R_R(R29) ,.T_L(T27), .T_R(T29), .R_old(R_old), .Z(Z28), .R(R28), .T(T28));
medianFilterCell  m29(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z28), .R_L(R28),.R_R(R30) ,.T_L(T28), .T_R(T30), .R_old(R_old), .Z(Z29), .R(R29), .T(T29));
medianFilterCell  m30(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z29), .R_L(R29),.R_R(R31) ,.T_L(T29), .T_R(T31), .R_old(R_old), .Z(Z30), .R(R30), .T(T30));
medianFilterCell  m31(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z30), .R_L(R30),.R_R(R32) ,.T_L(T30), .T_R(T32), .R_old(R_old), .Z(Z31), .R(R31), .T(T31));
medianFilterCell  m32(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z31), .R_L(R31),.R_R(R33) ,.T_L(T31), .T_R(T33), .R_old(R_old), .Z(Z32), .R(R32), .T(T32));
medianFilterCell  m33(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z32), .R_L(R32),.R_R(R34) ,.T_L(T32), .T_R(T34), .R_old(R_old), .Z(Z33), .R(R33), .T(T33));
medianFilterCell  m34(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z33), .R_L(R33),.R_R(R35) ,.T_L(T33), .T_R(T35), .R_old(R_old), .Z(Z34), .R(R34), .T(T34));
medianFilterCell  m35(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z34), .R_L(R34),.R_R(R36) ,.T_L(T34), .T_R(T36), .R_old(R_old), .Z(Z35), .R(R35), .T(T35));
medianFilterCell  m36(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z35), .R_L(R35),.R_R(R37) ,.T_L(T35), .T_R(T37), .R_old(R_old), .Z(Z36), .R(R36), .T(T36));
medianFilterCell  m37(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z36), .R_L(R36),.R_R(R38) ,.T_L(T36), .T_R(T38), .R_old(R_old), .Z(Z37), .R(R37), .T(T37));
medianFilterCell  m38(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z37), .R_L(R37),.R_R(R39) ,.T_L(T37), .T_R(T39), .R_old(R_old), .Z(Z38), .R(R38), .T(T38));
medianFilterCell  m39(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z38), .R_L(R38),.R_R(R40) ,.T_L(T38), .T_R(T40), .R_old(R_old), .Z(Z39), .R(R39), .T(T39));
medianFilterCell  m40(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z39), .R_L(R39),.R_R(R41) ,.T_L(T39), .T_R(T41), .R_old(R_old), .Z(Z40), .R(R40), .T(T40));
medianFilterCell  m41(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z40), .R_L(R40),.R_R(R42) ,.T_L(T40), .T_R(T42), .R_old(R_old), .Z(Z41), .R(R41), .T(T41));
medianFilterCell  m42(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z41), .R_L(R41),.R_R(R43) ,.T_L(T41), .T_R(T43), .R_old(R_old), .Z(Z42), .R(R42), .T(T42));
medianFilterCell  m43(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z42), .R_L(R42),.R_R(R44) ,.T_L(T42), .T_R(T44), .R_old(R_old), .Z(Z43), .R(R43), .T(T43));
medianFilterCell  m44(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z43), .R_L(R43),.R_R(R45) ,.T_L(T43), .T_R(T45), .R_old(R_old), .Z(Z44), .R(R44), .T(T44));
medianFilterCell  m45(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z44), .R_L(R44),.R_R(R46) ,.T_L(T44), .T_R(T46), .R_old(R_old), .Z(Z45), .R(R45), .T(T45));
medianFilterCell  m46(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z45), .R_L(R45),.R_R(R47) ,.T_L(T45), .T_R(T47), .R_old(R_old), .Z(Z46), .R(R46), .T(T46));
medianFilterCell  m47(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z46), .R_L(R46),.R_R(R48) ,.T_L(T46), .T_R(T48), .R_old(R_old), .Z(Z47), .R(R47), .T(T47));
medianFilterCell  m48(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z47), .R_L(R47),.R_R(R49) ,.T_L(T47), .T_R(T49), .R_old(R_old), .Z(Z48), .R(R48), .T(T48));
medianFilterCell  m49(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z48), .R_L(R48),.R_R(R50) ,.T_L(T48), .T_R(T50), .R_old(R_old), .Z(Z49), .R(R49), .T(T49));
medianFilterCell  m50(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z49), .R_L(R49),.R_R(R51) ,.T_L(T49), .T_R(T51), .R_old(R_old), .Z(Z50), .R(R50), .T(T50));
medianFilterCell  m51(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z50), .R_L(R50),.R_R(R52) ,.T_L(T50), .T_R(T52), .R_old(R_old), .Z(Z51), .R(R51), .T(T51));
medianFilterCell  m52(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z51), .R_L(R51),.R_R(R53) ,.T_L(T51), .T_R(T53), .R_old(R_old), .Z(Z52), .R(R52), .T(T52));
medianFilterCell  m53(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z52), .R_L(R52),.R_R(R54) ,.T_L(T52), .T_R(T54), .R_old(R_old), .Z(Z53), .R(R53), .T(T53));
medianFilterCell  m54(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z53), .R_L(R53),.R_R(R55) ,.T_L(T53), .T_R(T55), .R_old(R_old), .Z(Z54), .R(R54), .T(T54));
medianFilterCell  m55(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z54), .R_L(R54),.R_R(R56) ,.T_L(T54), .T_R(T56), .R_old(R_old), .Z(Z55), .R(R55), .T(T55));
medianFilterCell  m56(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z55), .R_L(R55),.R_R(R57) ,.T_L(T55), .T_R(T57), .R_old(R_old), .Z(Z56), .R(R56), .T(T56));
medianFilterCell  m57(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z56), .R_L(R56),.R_R(R58) ,.T_L(T56), .T_R(T58), .R_old(R_old), .Z(Z57), .R(R57), .T(T57));
medianFilterCell  m58(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z57), .R_L(R57),.R_R(R59) ,.T_L(T57), .T_R(T59), .R_old(R_old), .Z(Z58), .R(R58), .T(T58));
medianFilterCell  m59(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z58), .R_L(R58),.R_R(R60) ,.T_L(T58), .T_R(T60), .R_old(R_old), .Z(Z59), .R(R59), .T(T59));
medianFilterCell  m60(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z59), .R_L(R59),.R_R(R61) ,.T_L(T59), .T_R(T61), .R_old(R_old), .Z(Z60), .R(R60), .T(T60));
medianFilterCell  m61(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z60), .R_L(R60),.R_R(R62) ,.T_L(T60), .T_R(T62), .R_old(R_old), .Z(Z61), .R(R61), .T(T61));
medianFilterCell  m62(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z61), .R_L(R61),.R_R(R63) ,.T_L(T61), .T_R(T63), .R_old(R_old), .Z(Z62), .R(R62), .T(T62));
medianFilterCell  m63(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z62), .R_L(R62),.R_R(R64) ,.T_L(T62), .T_R(T64), .R_old(R_old), .Z(Z63), .R(R63), .T(T63));
medianFilterCell  m64(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z63), .R_L(R63),.R_R(R65) ,.T_L(T63), .T_R(T65), .R_old(R_old), .Z(Z64), .R(R64), .T(T64));
medianFilterCell  m65(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z64), .R_L(R64),.R_R(R66) ,.T_L(T64), .T_R(T66), .R_old(R_old), .Z(Z65), .R(R65), .T(T65));
medianFilterCell  m66(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z65), .R_L(R65),.R_R(R67) ,.T_L(T65), .T_R(T67), .R_old(R_old), .Z(Z66), .R(R66), .T(T66));
medianFilterCell  m67(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z66), .R_L(R66),.R_R(R68) ,.T_L(T66), .T_R(T68), .R_old(R_old), .Z(Z67), .R(R67), .T(T67));
medianFilterCell  m68(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z67), .R_L(R67),.R_R(R69) ,.T_L(T67), .T_R(T69), .R_old(R_old), .Z(Z68), .R(R68), .T(T68));
medianFilterCell  m69(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z68), .R_L(R68),.R_R(R70) ,.T_L(T68), .T_R(T70), .R_old(R_old), .Z(Z69), .R(R69), .T(T69));
medianFilterCell  m70(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z69), .R_L(R69),.R_R(R71) ,.T_L(T69), .T_R(T71), .R_old(R_old), .Z(Z70), .R(R70), .T(T70));
medianFilterCell  m71(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z70), .R_L(R70),.R_R(R72) ,.T_L(T70), .T_R(T72), .R_old(R_old), .Z(Z71), .R(R71), .T(T71));
medianFilterCell  m72(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z71), .R_L(R71),.R_R(R73) ,.T_L(T71), .T_R(T73), .R_old(R_old), .Z(Z72), .R(R72), .T(T72));
medianFilterCell  m73(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z72), .R_L(R72),.R_R(R74) ,.T_L(T72), .T_R(T74), .R_old(R_old), .Z(Z73), .R(R73), .T(T73));
medianFilterCell  m74(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z73), .R_L(R73),.R_R(R75) ,.T_L(T73), .T_R(T75), .R_old(R_old), .Z(Z74), .R(R74), .T(T74));
medianFilterCell  m75(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z74), .R_L(R74),.R_R(R76) ,.T_L(T74), .T_R(T76), .R_old(R_old), .Z(Z75), .R(R75), .T(T75));
medianFilterCell  m76(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z75), .R_L(R75),.R_R(R77) ,.T_L(T75), .T_R(T77), .R_old(R_old), .Z(Z76), .R(R76), .T(T76));
medianFilterCell  m77(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z76), .R_L(R76),.R_R(R78) ,.T_L(T76), .T_R(T78), .R_old(R_old), .Z(Z77), .R(R77), .T(T77));
medianFilterCell  m78(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z77), .R_L(R77),.R_R(R79) ,.T_L(T77), .T_R(T79), .R_old(R_old), .Z(Z78), .R(R78), .T(T78));
medianFilterCell  m79(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z78), .R_L(R78),.R_R(R80) ,.T_L(T78), .T_R(T80), .R_old(R_old), .Z(Z79), .R(R79), .T(T79));
medianFilterCell  m80(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z79), .R_L(R79),.R_R(R81) ,.T_L(T79), .T_R(T81), .R_old(R_old), .Z(Z80), .R(R80), .T(T80));
medianFilterCell  m81(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z80), .R_L(R80),.R_R(R82) ,.T_L(T80), .T_R(T82), .R_old(R_old), .Z(Z81), .R(R81), .T(T81));
medianFilterCell  m82(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z81), .R_L(R81),.R_R(R83) ,.T_L(T81), .T_R(T83), .R_old(R_old), .Z(Z82), .R(R82), .T(T82));
medianFilterCell  m83(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z82), .R_L(R82),.R_R(R84) ,.T_L(T82), .T_R(T84), .R_old(R_old), .Z(Z83), .R(R83), .T(T83));
medianFilterCell  m84(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z83), .R_L(R83),.R_R(R85) ,.T_L(T83), .T_R(T85), .R_old(R_old), .Z(Z84), .R(R84), .T(T84));
medianFilterCell  m85(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z84), .R_L(R84),.R_R(R86) ,.T_L(T84), .T_R(T86), .R_old(R_old), .Z(Z85), .R(R85), .T(T85));
medianFilterCell  m86(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z85), .R_L(R85),.R_R(R87) ,.T_L(T85), .T_R(T87), .R_old(R_old), .Z(Z86), .R(R86), .T(T86));
medianFilterCell  m87(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z86), .R_L(R86),.R_R(R88) ,.T_L(T86), .T_R(T88), .R_old(R_old), .Z(Z87), .R(R87), .T(T87));
medianFilterCell  m88(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z87), .R_L(R87),.R_R(R89) ,.T_L(T87), .T_R(T89), .R_old(R_old), .Z(Z88), .R(R88), .T(T88));
medianFilterCell  m89(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z88), .R_L(R88),.R_R(R90) ,.T_L(T88), .T_R(T90), .R_old(R_old), .Z(Z89), .R(R89), .T(T89));
medianFilterCell  m90(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z89), .R_L(R89),.R_R(R91) ,.T_L(T89), .T_R(T91), .R_old(R_old), .Z(Z90), .R(R90), .T(T90));
medianFilterCell  m91(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z90), .R_L(R90),.R_R(R92) ,.T_L(T90), .T_R(T92), .R_old(R_old), .Z(Z91), .R(R91), .T(T91));
medianFilterCell  m92(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z91), .R_L(R91),.R_R(R93) ,.T_L(T91), .T_R(T93), .R_old(R_old), .Z(Z92), .R(R92), .T(T92));
medianFilterCell  m93(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z92), .R_L(R92),.R_R(R94) ,.T_L(T92), .T_R(T94), .R_old(R_old), .Z(Z93), .R(R93), .T(T93));
medianFilterCell  m94(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z93), .R_L(R93),.R_R(R95) ,.T_L(T93), .T_R(T95), .R_old(R_old), .Z(Z94), .R(R94), .T(T94));
medianFilterCell  m95(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z94), .R_L(R94),.R_R(R96) ,.T_L(T94), .T_R(T96), .R_old(R_old), .Z(Z95), .R(R95), .T(T95));
medianFilterCell  m96(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z95), .R_L(R95),.R_R(R97) ,.T_L(T95), .T_R(T97), .R_old(R_old), .Z(Z96), .R(R96), .T(T96));
medianFilterCell  m97(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z96), .R_L(R96),.R_R(R98) ,.T_L(T96), .T_R(T98), .R_old(R_old), .Z(Z97), .R(R97), .T(T97));
medianFilterCell  m98(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z97), .R_L(R97),.R_R(R99) ,.T_L(T97), .T_R(T99), .R_old(R_old), .Z(Z98), .R(R98), .T(T98));
medianFilterCell  m99(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z98), .R_L(R98),.R_R(R100) ,.T_L(T98), .T_R(T100), .R_old(R_old), .Z(Z99), .R(R99), .T(T99));
medianFilterCell  m100(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z99), .R_L(R99),.R_R(R101) ,.T_L(T99), .T_R(T101), .R_old(R_old), .Z(Z100), .R(R100), .T(T100));
medianFilterCell  m101(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z100), .R_L(R100),.R_R(R102) ,.T_L(T100), .T_R(T102), .R_old(R_old), .Z(Z101), .R(R101), .T(T101));
medianFilterCell  m102(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z101), .R_L(R101),.R_R(R103) ,.T_L(T101), .T_R(T103), .R_old(R_old), .Z(Z102), .R(R102), .T(T102));
medianFilterCell  m103(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z102), .R_L(R102),.R_R(R104) ,.T_L(T102), .T_R(T104), .R_old(R_old), .Z(Z103), .R(R103), .T(T103));
medianFilterCell  m104(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z103), .R_L(R103),.R_R(R105) ,.T_L(T103), .T_R(T105), .R_old(R_old), .Z(Z104), .R(R104), .T(T104));
medianFilterCell  m105(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z104), .R_L(R104),.R_R(R106) ,.T_L(T104), .T_R(T106), .R_old(R_old), .Z(Z105), .R(R105), .T(T105));
medianFilterCell  m106(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z105), .R_L(R105),.R_R(R107) ,.T_L(T105), .T_R(T107), .R_old(R_old), .Z(Z106), .R(R106), .T(T106));
medianFilterCell  m107(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z106), .R_L(R106),.R_R(R108) ,.T_L(T106), .T_R(T108), .R_old(R_old), .Z(Z107), .R(R107), .T(T107));
medianFilterCell  m108(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z107), .R_L(R107),.R_R(R109) ,.T_L(T107), .T_R(T109), .R_old(R_old), .Z(Z108), .R(R108), .T(T108));
medianFilterCell  m109(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z108), .R_L(R108),.R_R(R110) ,.T_L(T108), .T_R(T110), .R_old(R_old), .Z(Z109), .R(R109), .T(T109));
medianFilterCell  m110(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z109), .R_L(R109),.R_R(R111) ,.T_L(T109), .T_R(T111), .R_old(R_old), .Z(Z110), .R(R110), .T(T110));
medianFilterCell  m111(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z110), .R_L(R110),.R_R(R112) ,.T_L(T110), .T_R(T112), .R_old(R_old), .Z(Z111), .R(R111), .T(T111));
medianFilterCell  m112(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z111), .R_L(R111),.R_R(R113) ,.T_L(T111), .T_R(T113), .R_old(R_old), .Z(Z112), .R(R112), .T(T112));
medianFilterCell  m113(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z112), .R_L(R112),.R_R(R114) ,.T_L(T112), .T_R(T114), .R_old(R_old), .Z(Z113), .R(R113), .T(T113));
medianFilterCell  m114(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z113), .R_L(R113),.R_R(R115) ,.T_L(T113), .T_R(T115), .R_old(R_old), .Z(Z114), .R(R114), .T(T114));
medianFilterCell  m115(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z114), .R_L(R114),.R_R(R116) ,.T_L(T114), .T_R(T116), .R_old(R_old), .Z(Z115), .R(R115), .T(T115));
medianFilterCell  m116(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z115), .R_L(R115),.R_R(R117) ,.T_L(T115), .T_R(T117), .R_old(R_old), .Z(Z116), .R(R116), .T(T116));
medianFilterCell  m117(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z116), .R_L(R116),.R_R(R118) ,.T_L(T116), .T_R(T118), .R_old(R_old), .Z(Z117), .R(R117), .T(T117));
medianFilterCell  m118(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z117), .R_L(R117),.R_R(R119) ,.T_L(T117), .T_R(T119), .R_old(R_old), .Z(Z118), .R(R118), .T(T118));
medianFilterCell  m119(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z118), .R_L(R118),.R_R(R120) ,.T_L(T118), .T_R(T120), .R_old(R_old), .Z(Z119), .R(R119), .T(T119));
medianFilterCell  m120(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z119), .R_L(R119),.R_R(R121) ,.T_L(T119), .T_R(T121), .R_old(R_old), .Z(Z120), .R(R120), .T(T120));
medianFilterCell  m121(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z120), .R_L(R120),.R_R(R122) ,.T_L(T120), .T_R(T122), .R_old(R_old), .Z(Z121), .R(R121), .T(T121));
medianFilterCell  m122(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z121), .R_L(R121),.R_R(R123) ,.T_L(T121), .T_R(T123), .R_old(R_old), .Z(Z122), .R(R122), .T(T122));
medianFilterCell  m123(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z122), .R_L(R122),.R_R(R124) ,.T_L(T122), .T_R(T124), .R_old(R_old), .Z(Z123), .R(R123), .T(T123));
medianFilterCell  m124(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z123), .R_L(R123),.R_R(R125) ,.T_L(T123), .T_R(T125), .R_old(R_old), .Z(Z124), .R(R124), .T(T124));
medianFilterCell  m125(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z124), .R_L(R124),.R_R(R126) ,.T_L(T124), .T_R(T126), .R_old(R_old), .Z(Z125), .R(R125), .T(T125));
medianFilterCell  m126(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z125), .R_L(R125),.R_R(R127) ,.T_L(T125), .T_R(T127), .R_old(R_old), .Z(Z126), .R(R126), .T(T126));
medianFilterCell  m127(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z126), .R_L(R126),.R_R(R128) ,.T_L(T126), .T_R(T128), .R_old(R_old), .Z(Z127), .R(R127), .T(T127));
medianFilterCell  m128(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z127), .R_L(R127),.R_R(R129) ,.T_L(T127), .T_R(T129), .R_old(R_old), .Z(Z128), .R(R128), .T(T128));
medianFilterCell  m129(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z128), .R_L(R128),.R_R(R130) ,.T_L(T128), .T_R(T130), .R_old(R_old), .Z(Z129), .R(R129), .T(T129));
medianFilterCell  m130(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z129), .R_L(R129),.R_R(R131) ,.T_L(T129), .T_R(T131), .R_old(R_old), .Z(Z130), .R(R130), .T(T130));
medianFilterCell  m131(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z130), .R_L(R130),.R_R(R132) ,.T_L(T130), .T_R(T132), .R_old(R_old), .Z(Z131), .R(R131), .T(T131));
medianFilterCell  m132(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z131), .R_L(R131),.R_R(R133) ,.T_L(T131), .T_R(T133), .R_old(R_old), .Z(Z132), .R(R132), .T(T132));
medianFilterCell  m133(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z132), .R_L(R132),.R_R(R134) ,.T_L(T132), .T_R(T134), .R_old(R_old), .Z(Z133), .R(R133), .T(T133));
medianFilterCell  m134(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z133), .R_L(R133),.R_R(R135) ,.T_L(T133), .T_R(T135), .R_old(R_old), .Z(Z134), .R(R134), .T(T134));
medianFilterCell  m135(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z134), .R_L(R134),.R_R(R136) ,.T_L(T134), .T_R(T136), .R_old(R_old), .Z(Z135), .R(R135), .T(T135));
medianFilterCell  m136(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z135), .R_L(R135),.R_R(R137) ,.T_L(T135), .T_R(T137), .R_old(R_old), .Z(Z136), .R(R136), .T(T136));
medianFilterCell  m137(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z136), .R_L(R136),.R_R(R138) ,.T_L(T136), .T_R(T138), .R_old(R_old), .Z(Z137), .R(R137), .T(T137));
medianFilterCell  m138(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z137), .R_L(R137),.R_R(R139) ,.T_L(T137), .T_R(T139), .R_old(R_old), .Z(Z138), .R(R138), .T(T138));
medianFilterCell  m139(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z138), .R_L(R138),.R_R(R140) ,.T_L(T138), .T_R(T140), .R_old(R_old), .Z(Z139), .R(R139), .T(T139));
medianFilterCell  m140(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z139), .R_L(R139),.R_R(R141) ,.T_L(T139), .T_R(T141), .R_old(R_old), .Z(Z140), .R(R140), .T(T140));
medianFilterCell  m141(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z140), .R_L(R140),.R_R(R142) ,.T_L(T140), .T_R(T142), .R_old(R_old), .Z(Z141), .R(R141), .T(T141));
medianFilterCell  m142(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z141), .R_L(R141),.R_R(R143) ,.T_L(T141), .T_R(T143), .R_old(R_old), .Z(Z142), .R(R142), .T(T142));
medianFilterCell  m143(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z142), .R_L(R142),.R_R(R144) ,.T_L(T142), .T_R(T144), .R_old(R_old), .Z(Z143), .R(R143), .T(T143));
medianFilterCell  m144(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z143), .R_L(R143),.R_R(R145) ,.T_L(T143), .T_R(T145), .R_old(R_old), .Z(Z144), .R(R144), .T(T144));
medianFilterCell  m145(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z144), .R_L(R144),.R_R(R146) ,.T_L(T144), .T_R(T146), .R_old(R_old), .Z(Z145), .R(R145), .T(T145));
medianFilterCell  m146(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z145), .R_L(R145),.R_R(R147) ,.T_L(T145), .T_R(T147), .R_old(R_old), .Z(Z146), .R(R146), .T(T146));
medianFilterCell  m147(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z146), .R_L(R146),.R_R(R148) ,.T_L(T146), .T_R(T148), .R_old(R_old), .Z(Z147), .R(R147), .T(T147));
medianFilterCell  m148(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z147), .R_L(R147),.R_R(R149) ,.T_L(T147), .T_R(T149), .R_old(R_old), .Z(Z148), .R(R148), .T(T148));
medianFilterCell  m149(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z148), .R_L(R148),.R_R(R150) ,.T_L(T148), .T_R(T150), .R_old(R_old), .Z(Z149), .R(R149), .T(T149));
medianFilterCell  m150(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z149), .R_L(R149),.R_R(R151) ,.T_L(T149), .T_R(T151), .R_old(R_old), .Z(Z150), .R(R150), .T(T150));
medianFilterCell  m151(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z150), .R_L(R150),.R_R(R152) ,.T_L(T150), .T_R(T152), .R_old(R_old), .Z(Z151), .R(R151), .T(T151));
medianFilterCell  m152(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z151), .R_L(R151),.R_R(R153) ,.T_L(T151), .T_R(T153), .R_old(R_old), .Z(Z152), .R(R152), .T(T152));
medianFilterCell  m153(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z152), .R_L(R152),.R_R(R154) ,.T_L(T152), .T_R(T154), .R_old(R_old), .Z(Z153), .R(R153), .T(T153));
medianFilterCell  m154(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z153), .R_L(R153),.R_R(R155) ,.T_L(T153), .T_R(T155), .R_old(R_old), .Z(Z154), .R(R154), .T(T154));
medianFilterCell  m155(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z154), .R_L(R154),.R_R(R156) ,.T_L(T154), .T_R(T156), .R_old(R_old), .Z(Z155), .R(R155), .T(T155));
medianFilterCell  m156(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z155), .R_L(R155),.R_R(R157) ,.T_L(T155), .T_R(T157), .R_old(R_old), .Z(Z156), .R(R156), .T(T156));
medianFilterCell  m157(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z156), .R_L(R156),.R_R(R158) ,.T_L(T156), .T_R(T158), .R_old(R_old), .Z(Z157), .R(R157), .T(T157));
medianFilterCell  m158(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z157), .R_L(R157),.R_R(R159) ,.T_L(T157), .T_R(T159), .R_old(R_old), .Z(Z158), .R(R158), .T(T158));
medianFilterCell  m159(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z158), .R_L(R158),.R_R(R160) ,.T_L(T158), .T_R(T160), .R_old(R_old), .Z(Z159), .R(R159), .T(T159));
medianFilterCell  m160(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z159), .R_L(R159),.R_R(R161) ,.T_L(T159), .T_R(T161), .R_old(R_old), .Z(Z160), .R(R160), .T(T160));
medianFilterCell  m161(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z160), .R_L(R160),.R_R(R162) ,.T_L(T160), .T_R(T162), .R_old(R_old), .Z(Z161), .R(R161), .T(T161));
medianFilterCell  m162(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z161), .R_L(R161),.R_R(R163) ,.T_L(T161), .T_R(T163), .R_old(R_old), .Z(Z162), .R(R162), .T(T162));
medianFilterCell  m163(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z162), .R_L(R162),.R_R(R164) ,.T_L(T162), .T_R(T164), .R_old(R_old), .Z(Z163), .R(R163), .T(T163));
medianFilterCell  m164(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z163), .R_L(R163),.R_R(R165) ,.T_L(T163), .T_R(T165), .R_old(R_old), .Z(Z164), .R(R164), .T(T164));
medianFilterCell  m165(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z164), .R_L(R164),.R_R(R166) ,.T_L(T164), .T_R(T166), .R_old(R_old), .Z(Z165), .R(R165), .T(T165));
medianFilterCell  m166(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z165), .R_L(R165),.R_R(R167) ,.T_L(T165), .T_R(T167), .R_old(R_old), .Z(Z166), .R(R166), .T(T166));
medianFilterCell  m167(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z166), .R_L(R166),.R_R(R168) ,.T_L(T166), .T_R(T168), .R_old(R_old), .Z(Z167), .R(R167), .T(T167));
medianFilterCell  m168(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z167), .R_L(R167),.R_R(R169) ,.T_L(T167), .T_R(T169), .R_old(R_old), .Z(Z168), .R(R168), .T(T168));
medianFilterCell  m169(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z168), .R_L(R168),.R_R(R170) ,.T_L(T168), .T_R(T170), .R_old(R_old), .Z(Z169), .R(R169), .T(T169));
medianFilterCell  m170(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z169), .R_L(R169),.R_R(R171) ,.T_L(T169), .T_R(T171), .R_old(R_old), .Z(Z170), .R(R170), .T(T170));
medianFilterCell  m171(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z170), .R_L(R170),.R_R(R172) ,.T_L(T170), .T_R(T172), .R_old(R_old), .Z(Z171), .R(R171), .T(T171));
medianFilterCell  m172(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z171), .R_L(R171),.R_R(R173) ,.T_L(T171), .T_R(T173), .R_old(R_old), .Z(Z172), .R(R172), .T(T172));
medianFilterCell  m173(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z172), .R_L(R172),.R_R(R174) ,.T_L(T172), .T_R(T174), .R_old(R_old), .Z(Z173), .R(R173), .T(T173));
medianFilterCell  m174(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z173), .R_L(R173),.R_R(R175) ,.T_L(T173), .T_R(T175), .R_old(R_old), .Z(Z174), .R(R174), .T(T174));
medianFilterCell  m175(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z174), .R_L(R174),.R_R(R176) ,.T_L(T174), .T_R(T176), .R_old(R_old), .Z(Z175), .R(R175), .T(T175));
medianFilterCell  m176(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z175), .R_L(R175),.R_R(R177) ,.T_L(T175), .T_R(T177), .R_old(R_old), .Z(Z176), .R(R176), .T(T176));
medianFilterCell  m177(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z176), .R_L(R176),.R_R(R178) ,.T_L(T176), .T_R(T178), .R_old(R_old), .Z(Z177), .R(R177), .T(T177));
medianFilterCell  m178(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z177), .R_L(R177),.R_R(R179) ,.T_L(T177), .T_R(T179), .R_old(R_old), .Z(Z178), .R(R178), .T(T178));
medianFilterCell  m179(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z178), .R_L(R178),.R_R(R180) ,.T_L(T178), .T_R(T180), .R_old(R_old), .Z(Z179), .R(R179), .T(T179));
medianFilterCell  m180(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z179), .R_L(R179),.R_R(R181) ,.T_L(T179), .T_R(T181), .R_old(R_old), .Z(Z180), .R(R180), .T(T180));
medianFilterCell  m181(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z180), .R_L(R180),.R_R(R182) ,.T_L(T180), .T_R(T182), .R_old(R_old), .Z(Z181), .R(R181), .T(T181));
medianFilterCell  m182(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z181), .R_L(R181),.R_R(R183) ,.T_L(T181), .T_R(T183), .R_old(R_old), .Z(Z182), .R(R182), .T(T182));
medianFilterCell  m183(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z182), .R_L(R182),.R_R(R184) ,.T_L(T182), .T_R(T184), .R_old(R_old), .Z(Z183), .R(R183), .T(T183));
medianFilterCell  m184(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z183), .R_L(R183),.R_R(R185) ,.T_L(T183), .T_R(T185), .R_old(R_old), .Z(Z184), .R(R184), .T(T184));
medianFilterCell  m185(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z184), .R_L(R184),.R_R(R186) ,.T_L(T184), .T_R(T186), .R_old(R_old), .Z(Z185), .R(R185), .T(T185));
medianFilterCell  m186(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z185), .R_L(R185),.R_R(R187) ,.T_L(T185), .T_R(T187), .R_old(R_old), .Z(Z186), .R(R186), .T(T186));
medianFilterCell  m187(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z186), .R_L(R186),.R_R(R188) ,.T_L(T186), .T_R(T188), .R_old(R_old), .Z(Z187), .R(R187), .T(T187));
medianFilterCell  m188(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z187), .R_L(R187),.R_R(R189) ,.T_L(T187), .T_R(T189), .R_old(R_old), .Z(Z188), .R(R188), .T(T188));
medianFilterCell  m189(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z188), .R_L(R188),.R_R(R190) ,.T_L(T188), .T_R(T190), .R_old(R_old), .Z(Z189), .R(R189), .T(T189));
medianFilterCell  m190(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z189), .R_L(R189),.R_R(R191) ,.T_L(T189), .T_R(T191), .R_old(R_old), .Z(Z190), .R(R190), .T(T190));
medianFilterCell  m191(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z190), .R_L(R190),.R_R(R192) ,.T_L(T190), .T_R(T192), .R_old(R_old), .Z(Z191), .R(R191), .T(T191));
medianFilterCell  m192(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z191), .R_L(R191),.R_R(R193) ,.T_L(T191), .T_R(T193), .R_old(R_old), .Z(Z192), .R(R192), .T(T192));
medianFilterCell  m193(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z192), .R_L(R192),.R_R(R194) ,.T_L(T192), .T_R(T194), .R_old(R_old), .Z(Z193), .R(R193), .T(T193));
medianFilterCell  m194(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z193), .R_L(R193),.R_R(R195) ,.T_L(T193), .T_R(T195), .R_old(R_old), .Z(Z194), .R(R194), .T(T194));
medianFilterCell  m195(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z194), .R_L(R194),.R_R(R196) ,.T_L(T194), .T_R(T196), .R_old(R_old), .Z(Z195), .R(R195), .T(T195));
medianFilterCell  m196(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z195), .R_L(R195),.R_R(R197) ,.T_L(T195), .T_R(T197), .R_old(R_old), .Z(Z196), .R(R196), .T(T196));
medianFilterCell  m197(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z196), .R_L(R196),.R_R(R198) ,.T_L(T196), .T_R(T198), .R_old(R_old), .Z(Z197), .R(R197), .T(T197));
medianFilterCell  m198(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z197), .R_L(R197),.R_R(R199) ,.T_L(T197), .T_R(T199), .R_old(R_old), .Z(Z198), .R(R198), .T(T198));
medianFilterCell  m199(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z198), .R_L(R198),.R_R(R200) ,.T_L(T198), .T_R(T200), .R_old(R_old), .Z(Z199), .R(R199), .T(T199));
medianFilterCell  m200(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z199), .R_L(R199),.R_R(R201) ,.T_L(T199), .T_R(T201), .R_old(R_old), .Z(Z200), .R(R200), .T(T200));
medianFilterCell  m201(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z200), .R_L(R200),.R_R(R202) ,.T_L(T200), .T_R(T202), .R_old(R_old), .Z(Z201), .R(R201), .T(T201));
medianFilterCell  m202(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z201), .R_L(R201),.R_R(R203) ,.T_L(T201), .T_R(T203), .R_old(R_old), .Z(Z202), .R(R202), .T(T202));
medianFilterCell  m203(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z202), .R_L(R202),.R_R(R204) ,.T_L(T202), .T_R(T204), .R_old(R_old), .Z(Z203), .R(R203), .T(T203));
medianFilterCell  m204(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z203), .R_L(R203),.R_R(R205) ,.T_L(T203), .T_R(T205), .R_old(R_old), .Z(Z204), .R(R204), .T(T204));
medianFilterCell  m205(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z204), .R_L(R204),.R_R(R206) ,.T_L(T204), .T_R(T206), .R_old(R_old), .Z(Z205), .R(R205), .T(T205));
medianFilterCell  m206(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z205), .R_L(R205),.R_R(R207) ,.T_L(T205), .T_R(T207), .R_old(R_old), .Z(Z206), .R(R206), .T(T206));
medianFilterCell  m207(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z206), .R_L(R206),.R_R(R208) ,.T_L(T206), .T_R(T208), .R_old(R_old), .Z(Z207), .R(R207), .T(T207));
medianFilterCell  m208(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z207), .R_L(R207),.R_R(R209) ,.T_L(T207), .T_R(T209), .R_old(R_old), .Z(Z208), .R(R208), .T(T208));
medianFilterCell  m209(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z208), .R_L(R208),.R_R(R210) ,.T_L(T208), .T_R(T210), .R_old(R_old), .Z(Z209), .R(R209), .T(T209));
medianFilterCell  m210(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z209), .R_L(R209),.R_R(R211) ,.T_L(T209), .T_R(T211), .R_old(R_old), .Z(Z210), .R(R210), .T(T210));
medianFilterCell  m211(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z210), .R_L(R210),.R_R(R212) ,.T_L(T210), .T_R(T212), .R_old(R_old), .Z(Z211), .R(R211), .T(T211));
medianFilterCell  m212(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z211), .R_L(R211),.R_R(R213) ,.T_L(T211), .T_R(T213), .R_old(R_old), .Z(Z212), .R(R212), .T(T212));
medianFilterCell  m213(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z212), .R_L(R212),.R_R(R214) ,.T_L(T212), .T_R(T214), .R_old(R_old), .Z(Z213), .R(R213), .T(T213));
medianFilterCell  m214(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z213), .R_L(R213),.R_R(R215) ,.T_L(T213), .T_R(T215), .R_old(R_old), .Z(Z214), .R(R214), .T(T214));
medianFilterCell  m215(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z214), .R_L(R214),.R_R(R216) ,.T_L(T214), .T_R(T216), .R_old(R_old), .Z(Z215), .R(R215), .T(T215));
medianFilterCell  m216(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z215), .R_L(R215),.R_R(R217) ,.T_L(T215), .T_R(T217), .R_old(R_old), .Z(Z216), .R(R216), .T(T216));
medianFilterCell  m217(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z216), .R_L(R216),.R_R(R218) ,.T_L(T216), .T_R(T218), .R_old(R_old), .Z(Z217), .R(R217), .T(T217));
medianFilterCell  m218(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z217), .R_L(R217),.R_R(R219) ,.T_L(T217), .T_R(T219), .R_old(R_old), .Z(Z218), .R(R218), .T(T218));
medianFilterCell  m219(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z218), .R_L(R218),.R_R(R220) ,.T_L(T218), .T_R(T220), .R_old(R_old), .Z(Z219), .R(R219), .T(T219));
medianFilterCell  m220(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z219), .R_L(R219),.R_R(R221) ,.T_L(T219), .T_R(T221), .R_old(R_old), .Z(Z220), .R(R220), .T(T220));
medianFilterCell  m221(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z220), .R_L(R220),.R_R(R222) ,.T_L(T220), .T_R(T222), .R_old(R_old), .Z(Z221), .R(R221), .T(T221));
medianFilterCell  m222(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z221), .R_L(R221),.R_R(R223) ,.T_L(T221), .T_R(T223), .R_old(R_old), .Z(Z222), .R(R222), .T(T222));
medianFilterCell  m223(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z222), .R_L(R222),.R_R(R224) ,.T_L(T222), .T_R(T224), .R_old(R_old), .Z(Z223), .R(R223), .T(T223));
medianFilterCell  m224(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z223), .R_L(R223),.R_R(R225) ,.T_L(T223), .T_R(T225), .R_old(R_old), .Z(Z224), .R(R224), .T(T224));
medianFilterCell  m225(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z224), .R_L(R224),.R_R(R226) ,.T_L(T224), .T_R(T226), .R_old(R_old), .Z(Z225), .R(R225), .T(T225));
medianFilterCell  m226(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z225), .R_L(R225),.R_R(R227) ,.T_L(T225), .T_R(T227), .R_old(R_old), .Z(Z226), .R(R226), .T(T226));
medianFilterCell  m227(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z226), .R_L(R226),.R_R(R228) ,.T_L(T226), .T_R(T228), .R_old(R_old), .Z(Z227), .R(R227), .T(T227));
medianFilterCell  m228(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z227), .R_L(R227),.R_R(R229) ,.T_L(T227), .T_R(T229), .R_old(R_old), .Z(Z228), .R(R228), .T(T228));
medianFilterCell  m229(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z228), .R_L(R228),.R_R(R230) ,.T_L(T228), .T_R(T230), .R_old(R_old), .Z(Z229), .R(R229), .T(T229));
medianFilterCell  m230(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z229), .R_L(R229),.R_R(R231) ,.T_L(T229), .T_R(T231), .R_old(R_old), .Z(Z230), .R(R230), .T(T230));
medianFilterCell  m231(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z230), .R_L(R230),.R_R(R232) ,.T_L(T230), .T_R(T232), .R_old(R_old), .Z(Z231), .R(R231), .T(T231));
medianFilterCell  m232(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z231), .R_L(R231),.R_R(R233) ,.T_L(T231), .T_R(T233), .R_old(R_old), .Z(Z232), .R(R232), .T(T232));
medianFilterCell  m233(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z232), .R_L(R232),.R_R(R234) ,.T_L(T232), .T_R(T234), .R_old(R_old), .Z(Z233), .R(R233), .T(T233));
medianFilterCell  m234(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z233), .R_L(R233),.R_R(R235) ,.T_L(T233), .T_R(T235), .R_old(R_old), .Z(Z234), .R(R234), .T(T234));
medianFilterCell  m235(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z234), .R_L(R234),.R_R(R236) ,.T_L(T234), .T_R(T236), .R_old(R_old), .Z(Z235), .R(R235), .T(T235));
medianFilterCell  m236(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z235), .R_L(R235),.R_R(R237) ,.T_L(T235), .T_R(T237), .R_old(R_old), .Z(Z236), .R(R236), .T(T236));
medianFilterCell  m237(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z236), .R_L(R236),.R_R(R238) ,.T_L(T236), .T_R(T238), .R_old(R_old), .Z(Z237), .R(R237), .T(T237));
medianFilterCell  m238(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z237), .R_L(R237),.R_R(R239) ,.T_L(T237), .T_R(T239), .R_old(R_old), .Z(Z238), .R(R238), .T(T238));
medianFilterCell  m239(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z238), .R_L(R238),.R_R(R240) ,.T_L(T238), .T_R(T240), .R_old(R_old), .Z(Z239), .R(R239), .T(T239));
medianFilterCell  m240(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z239), .R_L(R239),.R_R(R241) ,.T_L(T239), .T_R(T241), .R_old(R_old), .Z(Z240), .R(R240), .T(T240));
medianFilterCell  m241(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z240), .R_L(R240),.R_R(R242) ,.T_L(T240), .T_R(T242), .R_old(R_old), .Z(Z241), .R(R241), .T(T241));
medianFilterCell  m242(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z241), .R_L(R241),.R_R(R243) ,.T_L(T241), .T_R(T243), .R_old(R_old), .Z(Z242), .R(R242), .T(T242));
medianFilterCell  m243(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z242), .R_L(R242),.R_R(R244) ,.T_L(T242), .T_R(T244), .R_old(R_old), .Z(Z243), .R(R243), .T(T243));
medianFilterCell  m244(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z243), .R_L(R243),.R_R(R245) ,.T_L(T243), .T_R(T245), .R_old(R_old), .Z(Z244), .R(R244), .T(T244));
medianFilterCell  m245(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z244), .R_L(R244),.R_R(R246) ,.T_L(T244), .T_R(T246), .R_old(R_old), .Z(Z245), .R(R245), .T(T245));
medianFilterCell  m246(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z245), .R_L(R245),.R_R(R247) ,.T_L(T245), .T_R(T247), .R_old(R_old), .Z(Z246), .R(R246), .T(T246));
medianFilterCell  m247(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z246), .R_L(R246),.R_R(R248) ,.T_L(T246), .T_R(T248), .R_old(R_old), .Z(Z247), .R(R247), .T(T247));
medianFilterCell  m248(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z247), .R_L(R247),.R_R(R249) ,.T_L(T247), .T_R(T249), .R_old(R_old), .Z(Z248), .R(R248), .T(T248));
medianFilterCell  m249(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z248), .R_L(R248),.R_R(R250) ,.T_L(T248), .T_R(T250), .R_old(R_old), .Z(Z249), .R(R249), .T(T249));
medianFilterCell  m250(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z249), .R_L(R249),.R_R(R251) ,.T_L(T249), .T_R(T251), .R_old(R_old), .Z(Z250), .R(R250), .T(T250));
medianFilterCell  m251(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z250), .R_L(R250),.R_R(R252) ,.T_L(T250), .T_R(T252), .R_old(R_old), .Z(Z251), .R(R251), .T(T251));
medianFilterCell  m252(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z251), .R_L(R251),.R_R(R253) ,.T_L(T251), .T_R(T253), .R_old(R_old), .Z(Z252), .R(R252), .T(T252));
medianFilterCell  m253(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z252), .R_L(R252),.R_R(R254) ,.T_L(T252), .T_R(T254), .R_old(R_old), .Z(Z253), .R(R253), .T(T253));
medianFilterCell  m254(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z253), .R_L(R253),.R_R(R255) ,.T_L(T253), .T_R(T255), .R_old(R_old), .Z(Z254), .R(R254), .T(T254));
medianFilterCell  m255(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z254), .R_L(R254),.R_R(R256) ,.T_L(T254), .T_R(T256), .R_old(R_old), .Z(Z255), .R(R255), .T(T255));
medianFilterCell  m256(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z255), .R_L(R255),.R_R(R257) ,.T_L(T255), .T_R(T257), .R_old(R_old), .Z(Z256), .R(R256), .T(T256));
medianFilterCell  m257(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z256), .R_L(R256),.R_R(R258) ,.T_L(T256), .T_R(T258), .R_old(R_old), .Z(Z257), .R(R257), .T(T257));
medianFilterCell  m258(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z257), .R_L(R257),.R_R(R259) ,.T_L(T257), .T_R(T259), .R_old(R_old), .Z(Z258), .R(R258), .T(T258));
medianFilterCell  m259(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z258), .R_L(R258),.R_R(R260) ,.T_L(T258), .T_R(T260), .R_old(R_old), .Z(Z259), .R(R259), .T(T259));
medianFilterCell  m260(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z259), .R_L(R259),.R_R(R261) ,.T_L(T259), .T_R(T261), .R_old(R_old), .Z(Z260), .R(R260), .T(T260));
medianFilterCell  m261(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z260), .R_L(R260),.R_R(R262) ,.T_L(T260), .T_R(T262), .R_old(R_old), .Z(Z261), .R(R261), .T(T261));
medianFilterCell  m262(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z261), .R_L(R261),.R_R(R263) ,.T_L(T261), .T_R(T263), .R_old(R_old), .Z(Z262), .R(R262), .T(T262));
medianFilterCell  m263(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z262), .R_L(R262),.R_R(R264) ,.T_L(T262), .T_R(T264), .R_old(R_old), .Z(Z263), .R(R263), .T(T263));
medianFilterCell  m264(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z263), .R_L(R263),.R_R(R265) ,.T_L(T263), .T_R(T265), .R_old(R_old), .Z(Z264), .R(R264), .T(T264));
medianFilterCell  m265(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z264), .R_L(R264),.R_R(R266) ,.T_L(T264), .T_R(T266), .R_old(R_old), .Z(Z265), .R(R265), .T(T265));
medianFilterCell  m266(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z265), .R_L(R265),.R_R(R267) ,.T_L(T265), .T_R(T267), .R_old(R_old), .Z(Z266), .R(R266), .T(T266));
medianFilterCell  m267(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z266), .R_L(R266),.R_R(R268) ,.T_L(T266), .T_R(T268), .R_old(R_old), .Z(Z267), .R(R267), .T(T267));
medianFilterCell  m268(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z267), .R_L(R267),.R_R(R269) ,.T_L(T267), .T_R(T269), .R_old(R_old), .Z(Z268), .R(R268), .T(T268));
medianFilterCell  m269(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z268), .R_L(R268),.R_R(R270) ,.T_L(T268), .T_R(T270), .R_old(R_old), .Z(Z269), .R(R269), .T(T269));
medianFilterCell  m270(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z269), .R_L(R269),.R_R(R271) ,.T_L(T269), .T_R(T271), .R_old(R_old), .Z(Z270), .R(R270), .T(T270));
medianFilterCell  m271(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z270), .R_L(R270),.R_R(R272) ,.T_L(T270), .T_R(T272), .R_old(R_old), .Z(Z271), .R(R271), .T(T271));
medianFilterCell  m272(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z271), .R_L(R271),.R_R(R273) ,.T_L(T271), .T_R(T273), .R_old(R_old), .Z(Z272), .R(R272), .T(T272));
medianFilterCell  m273(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z272), .R_L(R272),.R_R(R274) ,.T_L(T272), .T_R(T274), .R_old(R_old), .Z(Z273), .R(R273), .T(T273));
medianFilterCell  m274(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z273), .R_L(R273),.R_R(R275) ,.T_L(T273), .T_R(T275), .R_old(R_old), .Z(Z274), .R(R274), .T(T274));
medianFilterCell  m275(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z274), .R_L(R274),.R_R(R276) ,.T_L(T274), .T_R(T276), .R_old(R_old), .Z(Z275), .R(R275), .T(T275));
medianFilterCell  m276(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z275), .R_L(R275),.R_R(R277) ,.T_L(T275), .T_R(T277), .R_old(R_old), .Z(Z276), .R(R276), .T(T276));
medianFilterCell  m277(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z276), .R_L(R276),.R_R(R278) ,.T_L(T276), .T_R(T278), .R_old(R_old), .Z(Z277), .R(R277), .T(T277));
medianFilterCell  m278(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z277), .R_L(R277),.R_R(R279) ,.T_L(T277), .T_R(T279), .R_old(R_old), .Z(Z278), .R(R278), .T(T278));
medianFilterCell  m279(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z278), .R_L(R278),.R_R(R280) ,.T_L(T278), .T_R(T280), .R_old(R_old), .Z(Z279), .R(R279), .T(T279));
medianFilterCell  m280(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z279), .R_L(R279),.R_R(R281) ,.T_L(T279), .T_R(T281), .R_old(R_old), .Z(Z280), .R(R280), .T(T280));
medianFilterCell  m281(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z280), .R_L(R280),.R_R(R282) ,.T_L(T280), .T_R(T282), .R_old(R_old), .Z(Z281), .R(R281), .T(T281));
medianFilterCell  m282(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z281), .R_L(R281),.R_R(R283) ,.T_L(T281), .T_R(T283), .R_old(R_old), .Z(Z282), .R(R282), .T(T282));
medianFilterCell  m283(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z282), .R_L(R282),.R_R(R284) ,.T_L(T282), .T_R(T284), .R_old(R_old), .Z(Z283), .R(R283), .T(T283));
medianFilterCell  m284(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z283), .R_L(R283),.R_R(R285) ,.T_L(T283), .T_R(T285), .R_old(R_old), .Z(Z284), .R(R284), .T(T284));
medianFilterCell  m285(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z284), .R_L(R284),.R_R(R286) ,.T_L(T284), .T_R(T286), .R_old(R_old), .Z(Z285), .R(R285), .T(T285));
medianFilterCell  m286(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z285), .R_L(R285),.R_R(R287) ,.T_L(T285), .T_R(T287), .R_old(R_old), .Z(Z286), .R(R286), .T(T286));
medianFilterCell  m287(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z286), .R_L(R286),.R_R(R288) ,.T_L(T286), .T_R(T288), .R_old(R_old), .Z(Z287), .R(R287), .T(T287));
medianFilterCell  m288(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z287), .R_L(R287),.R_R(R289) ,.T_L(T287), .T_R(T289), .R_old(R_old), .Z(Z288), .R(R288), .T(T288));
medianFilterCell  m289(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z288), .R_L(R288),.R_R(R290) ,.T_L(T288), .T_R(T290), .R_old(R_old), .Z(Z289), .R(R289), .T(T289));
medianFilterCell  m290(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z289), .R_L(R289),.R_R(R291) ,.T_L(T289), .T_R(T291), .R_old(R_old), .Z(Z290), .R(R290), .T(T290));
medianFilterCell  m291(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z290), .R_L(R290),.R_R(R292) ,.T_L(T290), .T_R(T292), .R_old(R_old), .Z(Z291), .R(R291), .T(T291));
medianFilterCell  m292(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z291), .R_L(R291),.R_R(R293) ,.T_L(T291), .T_R(T293), .R_old(R_old), .Z(Z292), .R(R292), .T(T292));
medianFilterCell  m293(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z292), .R_L(R292),.R_R(R294) ,.T_L(T292), .T_R(T294), .R_old(R_old), .Z(Z293), .R(R293), .T(T293));
medianFilterCell  m294(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z293), .R_L(R293),.R_R(R295) ,.T_L(T293), .T_R(T295), .R_old(R_old), .Z(Z294), .R(R294), .T(T294));
medianFilterCell  m295(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z294), .R_L(R294),.R_R(R296) ,.T_L(T294), .T_R(T296), .R_old(R_old), .Z(Z295), .R(R295), .T(T295));
medianFilterCell  m296(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z295), .R_L(R295),.R_R(R297) ,.T_L(T295), .T_R(T297), .R_old(R_old), .Z(Z296), .R(R296), .T(T296));
medianFilterCell  m297(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z296), .R_L(R296),.R_R(R298) ,.T_L(T296), .T_R(T298), .R_old(R_old), .Z(Z297), .R(R297), .T(T297));
medianFilterCell  m298(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z297), .R_L(R297),.R_R(R299) ,.T_L(T297), .T_R(T299), .R_old(R_old), .Z(Z298), .R(R298), .T(T298));
medianFilterCell  m299(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z298), .R_L(R298),.R_R(R300) ,.T_L(T298), .T_R(T300), .R_old(R_old), .Z(Z299), .R(R299), .T(T299));
medianCell_rightMst  m300(.X(X) ,.clk(clk), .reset(reset), .Z_L(Z299), .R_L(R299), .T_L(T299), .R(R300),.T(T300));


endmodule