`ifndef _my_include_vh_
`define _my_include_vh_

