`timescale 1ns / 1ps
`include "macro.vh"
///////////////////////
module top ( clk ,reset ,X ,median );

output [`DATA_LENGTH-1:0] median ;
input [`DATA_LENGTH-1:0] X ;
input clk ,reset ;
reg  flag ;
reg [`DATA_LENGTH-1:0] median;wire  [`DATA_LENGTH-1:0] oldData ;
wire 	[`DATA_LENGTH-1:0] dataOut1 ,dataOut2 ,dataOut3 ,dataOut4 ,dataOut5 ,dataOut6 ,dataOut7 ,dataOut8 ,dataOut9 ,dataOut10 ,dataOut11 ,dataOut12 ,dataOut13 ,dataOut14 ,dataOut15 ,dataOut16 ,dataOut17 ,dataOut18 ,dataOut19 ,dataOut20 ,dataOut21 ,dataOut22 ,dataOut23 ,dataOut24 ,dataOut25 ,dataOut26 ,dataOut27 ,dataOut28 ,dataOut29 ,dataOut30 ,dataOut31 ,dataOut32 ,dataOut33 ,dataOut34 ,dataOut35 ,dataOut36 ,dataOut37 ,dataOut38 ,dataOut39 ,dataOut40 ,dataOut41 ,dataOut42 ,dataOut43 ,dataOut44 ,dataOut45 ,dataOut46 ,dataOut47 ,dataOut48 ,dataOut49 ,dataOut50 ,dataOut51 ,dataOut52 ,dataOut53 ,dataOut54 ,dataOut55 ,dataOut56 ,dataOut57 ,dataOut58 ,dataOut59 ,dataOut60 ,dataOut61 ,dataOut62 ,dataOut63 ,dataOut64 ,dataOut65 ,dataOut66 ,dataOut67 ,dataOut68 ,dataOut69 ,dataOut70 ,dataOut71 ,dataOut72 ,dataOut73 ,dataOut74 ,dataOut75 ,dataOut76 ,dataOut77 ,dataOut78 ,dataOut79 ,dataOut80 ,dataOut81 ,dataOut82 ,dataOut83 ,dataOut84 ,dataOut85 ,dataOut86 ,dataOut87 ,dataOut88 ,dataOut89 ,dataOut90 ,dataOut91 ,dataOut92 ,dataOut93 ,dataOut94 ,dataOut95 ,dataOut96 ,dataOut97 ,dataOut98 ,dataOut99 ,dataOut100 ,dataOut101 ,dataOut102 ,dataOut103 ,dataOut104 ,dataOut105 ,dataOut106 ,dataOut107 ,dataOut108 ,dataOut109 ,dataOut110 ,dataOut111 ,dataOut112 ,dataOut113 ,dataOut114 ,dataOut115 ,dataOut116 ,dataOut117 ,dataOut118 ,dataOut119 ,dataOut120 ,dataOut121 ,dataOut122 ,dataOut123 ,dataOut124 ,dataOut125 ,dataOut126 ,dataOut127 ,dataOut128 ,dataOut129 ,dataOut130 ,dataOut131 ,dataOut132 ,dataOut133 ,dataOut134 ,dataOut135 ,dataOut136 ,dataOut137 ,dataOut138 ,dataOut139 ,dataOut140 ,dataOut141 ,dataOut142 ,dataOut143 ,dataOut144 ,dataOut145 ,dataOut146 ,dataOut147 ,dataOut148 ,dataOut149 ,dataOut150 ,dataOut151 ,dataOut152 ,dataOut153 ,dataOut154 ,dataOut155 ,dataOut156 ,dataOut157 ,dataOut158 ,dataOut159 ,dataOut160 ,dataOut161 ,dataOut162 ,dataOut163 ,dataOut164 ,dataOut165 ,dataOut166 ,dataOut167 ,dataOut168 ,dataOut169 ,dataOut170 ,dataOut171 ,dataOut172 ,dataOut173 ,dataOut174 ,dataOut175 ,dataOut176 ,dataOut177 ,dataOut178 ,dataOut179 ,dataOut180 ,dataOut181 ,dataOut182 ,dataOut183 ,dataOut184 ,dataOut185 ,dataOut186 ,dataOut187 ,dataOut188 ,dataOut189 ,dataOut190 ,dataOut191 ,dataOut192 ,dataOut193 ,dataOut194 ,dataOut195 ,dataOut196 ,dataOut197 ,dataOut198 ,dataOut199 ,dataOut200 ,dataOut201 ,dataOut202 ,dataOut203 ,dataOut204 ,dataOut205 ,dataOut206 ,dataOut207 ,dataOut208 ,dataOut209 ,dataOut210 ,dataOut211 ,dataOut212 ,dataOut213 ,dataOut214 ,dataOut215 ,dataOut216 ,dataOut217 ,dataOut218 ,dataOut219 ,dataOut220 ,dataOut221 ,dataOut222 ,dataOut223 ,dataOut224 ,dataOut225 ,dataOut226 ,dataOut227 ,dataOut228 ,dataOut229 ,dataOut230 ,dataOut231 ,dataOut232 ,dataOut233 ,dataOut234 ,dataOut235 ,dataOut236 ,dataOut237 ,dataOut238 ,dataOut239 ,dataOut240 ,dataOut241 ,dataOut242 ,dataOut243 ,dataOut244 ,dataOut245 ,dataOut246 ,dataOut247 ,dataOut248 ,dataOut249 ,dataOut250 ,dataOut251 ,dataOut252 ,dataOut253 ,dataOut254 ,dataOut255 ,dataOut256 ,dataOut257 ,dataOut258 ,dataOut259 ,dataOut260 ,dataOut261 ,dataOut262 ,dataOut263 ,dataOut264 ,dataOut265 ,dataOut266 ,dataOut267 ,dataOut268 ,dataOut269 ,dataOut270 ,dataOut271 ,dataOut272 ,dataOut273 ,dataOut274 ,dataOut275 ,dataOut276 ,dataOut277 ,dataOut278 ,dataOut279 ,dataOut280 ,dataOut281 ,dataOut282 ,dataOut283 ,dataOut284 ,dataOut285 ,dataOut286 ,dataOut287 ,dataOut288 ,dataOut289 ,dataOut290 ,dataOut291 ,dataOut292 ,dataOut293 ,dataOut294 ,dataOut295 ,dataOut296 ,dataOut297 ,dataOut298 ,dataOut299 ,dataOut300 ,dataOut301 ,dataOut302 ,dataOut303 ,dataOut304 ,dataOut305 ,dataOut306 ,dataOut307 ,dataOut308 ,dataOut309 ,dataOut310 ,dataOut311 ,dataOut312 ,dataOut313 ,dataOut314 ,dataOut315 ,dataOut316 ,dataOut317 ,dataOut318 ,dataOut319 ,dataOut320 ,dataOut321 ,dataOut322 ,dataOut323 ,dataOut324 ,dataOut325 ,dataOut326 ,dataOut327 ,dataOut328 ,dataOut329 ,dataOut330 ,dataOut331 ,dataOut332 ,dataOut333 ,dataOut334 ,dataOut335 ,dataOut336 ,dataOut337 ,dataOut338 ,dataOut339 ,dataOut340 ,dataOut341 ,dataOut342 ,dataOut343 ,dataOut344 ,dataOut345 ,dataOut346 ,dataOut347 ,dataOut348 ,dataOut349 ,dataOut350 ,dataOut351 ,dataOut352 ,dataOut353 ,dataOut354 ,dataOut355 ,dataOut356 ,dataOut357 ,dataOut358 ,dataOut359 ,dataOut360 ,dataOut361 ,dataOut362 ,dataOut363 ,dataOut364 ,dataOut365 ,dataOut366 ,dataOut367 ,dataOut368 ,dataOut369 ,dataOut370 ,dataOut371 ,dataOut372 ,dataOut373 ,dataOut374 ,dataOut375 ,dataOut376 ,dataOut377 ,dataOut378 ,dataOut379 ,dataOut380 ,dataOut381 ,dataOut382 ,dataOut383 ,dataOut384 ,dataOut385 ,dataOut386 ,dataOut387 ,dataOut388 ,dataOut389 ,dataOut390 ,dataOut391 ,dataOut392 ,dataOut393 ,dataOut394 ,dataOut395 ,dataOut396 ,dataOut397 ,dataOut398 ,dataOut399 ,dataOut400 ,dataOut401 ,dataOut402 ,dataOut403 ,dataOut404 ,dataOut405 ,dataOut406 ,dataOut407 ,dataOut408 ,dataOut409 ,dataOut410 ,dataOut411 ,dataOut412 ,dataOut413 ,dataOut414 ,dataOut415 ,dataOut416 ,dataOut417 ,dataOut418 ,dataOut419 ,dataOut420 ,dataOut421 ,dataOut422 ,dataOut423 ,dataOut424 ,dataOut425 ,dataOut426 ,dataOut427 ,dataOut428 ,dataOut429 ,dataOut430 ,dataOut431 ,dataOut432 ,dataOut433 ,dataOut434 ,dataOut435 ,dataOut436 ,dataOut437 ,dataOut438 ,dataOut439 ,dataOut440 ,dataOut441 ,dataOut442 ,dataOut443 ,dataOut444 ,dataOut445 ,dataOut446 ,dataOut447 ,dataOut448 ,dataOut449 ,dataOut450 ,dataOut451 ,dataOut452 ,dataOut453 ,dataOut454 ,dataOut455 ,dataOut456 ,dataOut457 ,dataOut458 ,dataOut459 ,dataOut460 ,dataOut461 ,dataOut462 ,dataOut463 ,dataOut464 ,dataOut465 ,dataOut466 ,dataOut467 ,dataOut468 ,dataOut469 ,dataOut470 ,dataOut471 ,dataOut472 ,dataOut473 ,dataOut474 ,dataOut475 ,dataOut476 ,dataOut477 ,dataOut478 ,dataOut479 ,dataOut480 ,dataOut481 ,dataOut482 ,dataOut483 ,dataOut484 ,dataOut485 ,dataOut486 ,dataOut487 ,dataOut488 ,dataOut489 ,dataOut490 ,dataOut491 ,dataOut492 ,dataOut493 ,dataOut494 ,dataOut495 ,dataOut496 ,dataOut497 ,dataOut498 ,dataOut499 ,dataOut500 ,dataOut501 ,dataOut502 ,dataOut503 ,dataOut504 ,dataOut505 ,dataOut506 ,dataOut507 ,dataOut508 ,dataOut509 ,dataOut510 ,dataOut511 ,dataOut512 ,dataOut513 ,dataOut514 ,dataOut515 ,dataOut516 ,dataOut517 ,dataOut518 ,dataOut519 ,dataOut520 ,dataOut521 ,dataOut522 ,dataOut523 ,dataOut524 ,dataOut525 ,dataOut526 ,dataOut527 ,dataOut528 ,dataOut529 ,dataOut530 ,dataOut531 ,dataOut532 ,dataOut533 ,dataOut534 ,dataOut535 ,dataOut536 ,dataOut537 ,dataOut538 ,dataOut539 ,dataOut540 ,dataOut541 ,dataOut542 ,dataOut543 ,dataOut544 ,dataOut545 ,dataOut546 ,dataOut547 ,dataOut548 ,dataOut549 ,dataOut550 ,dataOut551 ,dataOut552 ,dataOut553 ,dataOut554 ,dataOut555 ,dataOut556 ,dataOut557 ,dataOut558 ,dataOut559 ,dataOut560 ,dataOut561 ,dataOut562 ,dataOut563 ,dataOut564 ,dataOut565 ,dataOut566 ,dataOut567 ,dataOut568 ,dataOut569 ,dataOut570 ,dataOut571 ,dataOut572 ,dataOut573 ,dataOut574 ,dataOut575 ,dataOut576 ,dataOut577 ,dataOut578 ,dataOut579 ,dataOut580 ,dataOut581 ,dataOut582 ,dataOut583 ,dataOut584 ,dataOut585 ,dataOut586 ,dataOut587 ,dataOut588 ,dataOut589 ,dataOut590 ,dataOut591 ,dataOut592 ,dataOut593 ,dataOut594 ,dataOut595 ,dataOut596 ,dataOut597 ,dataOut598 ,dataOut599 ,dataOut600 ,dataOut601 ,dataOut602 ,dataOut603 ,dataOut604 ,dataOut605 ,dataOut606 ,dataOut607 ,dataOut608 ,dataOut609 ,dataOut610 ,dataOut611 ,dataOut612 ,dataOut613 ,dataOut614 ,dataOut615 ,dataOut616 ,dataOut617 ,dataOut618 ,dataOut619 ,dataOut620 ,dataOut621 ,dataOut622 ,dataOut623 ,dataOut624 ,dataOut625 ,dataOut626 ,dataOut627 ,dataOut628 ,dataOut629 ,dataOut630 ,dataOut631 ,dataOut632 ,dataOut633 ,dataOut634 ,dataOut635 ,dataOut636 ,dataOut637 ,dataOut638 ,dataOut639 ,dataOut640 ,dataOut641 ,dataOut642 ,dataOut643 ,dataOut644 ,dataOut645 ,dataOut646 ,dataOut647 ,dataOut648 ,dataOut649 ,dataOut650 ,dataOut651 ,dataOut652 ,dataOut653 ,dataOut654 ,dataOut655 ,dataOut656 ,dataOut657 ,dataOut658 ,dataOut659 ,dataOut660 ,dataOut661 ,dataOut662 ,dataOut663 ,dataOut664 ,dataOut665 ,dataOut666 ,dataOut667 ,dataOut668 ,dataOut669 ,dataOut670 ,dataOut671 ,dataOut672 ,dataOut673 ,dataOut674 ,dataOut675 ,dataOut676 ,dataOut677 ,dataOut678 ,dataOut679 ,dataOut680 ,dataOut681 ,dataOut682 ,dataOut683 ,dataOut684 ,dataOut685 ,dataOut686 ,dataOut687 ,dataOut688 ,dataOut689 ,dataOut690 ,dataOut691 ,dataOut692 ,dataOut693 ,dataOut694 ,dataOut695 ,dataOut696 ,dataOut697 ,dataOut698 ,dataOut699 ,dataOut700;
wire 	 R1 ,R2 ,R3 ,R4 ,R5 ,R6 ,R7 ,R8 ,R9 ,R10 ,R11 ,R12 ,R13 ,R14 ,R15 ,R16 ,R17 ,R18 ,R19 ,R20 ,R21 ,R22 ,R23 ,R24 ,R25 ,R26 ,R27 ,R28 ,R29 ,R30 ,R31 ,R32 ,R33 ,R34 ,R35 ,R36 ,R37 ,R38 ,R39 ,R40 ,R41 ,R42 ,R43 ,R44 ,R45 ,R46 ,R47 ,R48 ,R49 ,R50 ,R51 ,R52 ,R53 ,R54 ,R55 ,R56 ,R57 ,R58 ,R59 ,R60 ,R61 ,R62 ,R63 ,R64 ,R65 ,R66 ,R67 ,R68 ,R69 ,R70 ,R71 ,R72 ,R73 ,R74 ,R75 ,R76 ,R77 ,R78 ,R79 ,R80 ,R81 ,R82 ,R83 ,R84 ,R85 ,R86 ,R87 ,R88 ,R89 ,R90 ,R91 ,R92 ,R93 ,R94 ,R95 ,R96 ,R97 ,R98 ,R99 ,R100 ,R101 ,R102 ,R103 ,R104 ,R105 ,R106 ,R107 ,R108 ,R109 ,R110 ,R111 ,R112 ,R113 ,R114 ,R115 ,R116 ,R117 ,R118 ,R119 ,R120 ,R121 ,R122 ,R123 ,R124 ,R125 ,R126 ,R127 ,R128 ,R129 ,R130 ,R131 ,R132 ,R133 ,R134 ,R135 ,R136 ,R137 ,R138 ,R139 ,R140 ,R141 ,R142 ,R143 ,R144 ,R145 ,R146 ,R147 ,R148 ,R149 ,R150 ,R151 ,R152 ,R153 ,R154 ,R155 ,R156 ,R157 ,R158 ,R159 ,R160 ,R161 ,R162 ,R163 ,R164 ,R165 ,R166 ,R167 ,R168 ,R169 ,R170 ,R171 ,R172 ,R173 ,R174 ,R175 ,R176 ,R177 ,R178 ,R179 ,R180 ,R181 ,R182 ,R183 ,R184 ,R185 ,R186 ,R187 ,R188 ,R189 ,R190 ,R191 ,R192 ,R193 ,R194 ,R195 ,R196 ,R197 ,R198 ,R199 ,R200 ,R201 ,R202 ,R203 ,R204 ,R205 ,R206 ,R207 ,R208 ,R209 ,R210 ,R211 ,R212 ,R213 ,R214 ,R215 ,R216 ,R217 ,R218 ,R219 ,R220 ,R221 ,R222 ,R223 ,R224 ,R225 ,R226 ,R227 ,R228 ,R229 ,R230 ,R231 ,R232 ,R233 ,R234 ,R235 ,R236 ,R237 ,R238 ,R239 ,R240 ,R241 ,R242 ,R243 ,R244 ,R245 ,R246 ,R247 ,R248 ,R249 ,R250 ,R251 ,R252 ,R253 ,R254 ,R255 ,R256 ,R257 ,R258 ,R259 ,R260 ,R261 ,R262 ,R263 ,R264 ,R265 ,R266 ,R267 ,R268 ,R269 ,R270 ,R271 ,R272 ,R273 ,R274 ,R275 ,R276 ,R277 ,R278 ,R279 ,R280 ,R281 ,R282 ,R283 ,R284 ,R285 ,R286 ,R287 ,R288 ,R289 ,R290 ,R291 ,R292 ,R293 ,R294 ,R295 ,R296 ,R297 ,R298 ,R299 ,R300 ,R301 ,R302 ,R303 ,R304 ,R305 ,R306 ,R307 ,R308 ,R309 ,R310 ,R311 ,R312 ,R313 ,R314 ,R315 ,R316 ,R317 ,R318 ,R319 ,R320 ,R321 ,R322 ,R323 ,R324 ,R325 ,R326 ,R327 ,R328 ,R329 ,R330 ,R331 ,R332 ,R333 ,R334 ,R335 ,R336 ,R337 ,R338 ,R339 ,R340 ,R341 ,R342 ,R343 ,R344 ,R345 ,R346 ,R347 ,R348 ,R349 ,R350 ,R351 ,R352 ,R353 ,R354 ,R355 ,R356 ,R357 ,R358 ,R359 ,R360 ,R361 ,R362 ,R363 ,R364 ,R365 ,R366 ,R367 ,R368 ,R369 ,R370 ,R371 ,R372 ,R373 ,R374 ,R375 ,R376 ,R377 ,R378 ,R379 ,R380 ,R381 ,R382 ,R383 ,R384 ,R385 ,R386 ,R387 ,R388 ,R389 ,R390 ,R391 ,R392 ,R393 ,R394 ,R395 ,R396 ,R397 ,R398 ,R399 ,R400 ,R401 ,R402 ,R403 ,R404 ,R405 ,R406 ,R407 ,R408 ,R409 ,R410 ,R411 ,R412 ,R413 ,R414 ,R415 ,R416 ,R417 ,R418 ,R419 ,R420 ,R421 ,R422 ,R423 ,R424 ,R425 ,R426 ,R427 ,R428 ,R429 ,R430 ,R431 ,R432 ,R433 ,R434 ,R435 ,R436 ,R437 ,R438 ,R439 ,R440 ,R441 ,R442 ,R443 ,R444 ,R445 ,R446 ,R447 ,R448 ,R449 ,R450 ,R451 ,R452 ,R453 ,R454 ,R455 ,R456 ,R457 ,R458 ,R459 ,R460 ,R461 ,R462 ,R463 ,R464 ,R465 ,R466 ,R467 ,R468 ,R469 ,R470 ,R471 ,R472 ,R473 ,R474 ,R475 ,R476 ,R477 ,R478 ,R479 ,R480 ,R481 ,R482 ,R483 ,R484 ,R485 ,R486 ,R487 ,R488 ,R489 ,R490 ,R491 ,R492 ,R493 ,R494 ,R495 ,R496 ,R497 ,R498 ,R499 ,R500 ,R501 ,R502 ,R503 ,R504 ,R505 ,R506 ,R507 ,R508 ,R509 ,R510 ,R511 ,R512 ,R513 ,R514 ,R515 ,R516 ,R517 ,R518 ,R519 ,R520 ,R521 ,R522 ,R523 ,R524 ,R525 ,R526 ,R527 ,R528 ,R529 ,R530 ,R531 ,R532 ,R533 ,R534 ,R535 ,R536 ,R537 ,R538 ,R539 ,R540 ,R541 ,R542 ,R543 ,R544 ,R545 ,R546 ,R547 ,R548 ,R549 ,R550 ,R551 ,R552 ,R553 ,R554 ,R555 ,R556 ,R557 ,R558 ,R559 ,R560 ,R561 ,R562 ,R563 ,R564 ,R565 ,R566 ,R567 ,R568 ,R569 ,R570 ,R571 ,R572 ,R573 ,R574 ,R575 ,R576 ,R577 ,R578 ,R579 ,R580 ,R581 ,R582 ,R583 ,R584 ,R585 ,R586 ,R587 ,R588 ,R589 ,R590 ,R591 ,R592 ,R593 ,R594 ,R595 ,R596 ,R597 ,R598 ,R599 ,R600 ,R601 ,R602 ,R603 ,R604 ,R605 ,R606 ,R607 ,R608 ,R609 ,R610 ,R611 ,R612 ,R613 ,R614 ,R615 ,R616 ,R617 ,R618 ,R619 ,R620 ,R621 ,R622 ,R623 ,R624 ,R625 ,R626 ,R627 ,R628 ,R629 ,R630 ,R631 ,R632 ,R633 ,R634 ,R635 ,R636 ,R637 ,R638 ,R639 ,R640 ,R641 ,R642 ,R643 ,R644 ,R645 ,R646 ,R647 ,R648 ,R649 ,R650 ,R651 ,R652 ,R653 ,R654 ,R655 ,R656 ,R657 ,R658 ,R659 ,R660 ,R661 ,R662 ,R663 ,R664 ,R665 ,R666 ,R667 ,R668 ,R669 ,R670 ,R671 ,R672 ,R673 ,R674 ,R675 ,R676 ,R677 ,R678 ,R679 ,R680 ,R681 ,R682 ,R683 ,R684 ,R685 ,R686 ,R687 ,R688 ,R689 ,R690 ,R691 ,R692 ,R693 ,R694 ,R695 ,R696 ,R697 ,R698 ,R699 ,R700;
always @(posedge clk or  posedge reset)
begin
	if(reset)
		flag <= 0;
	else
	begin
		flag <= ~flag ;
		if (flag ==0)
			 median <= (dataOut350 + dataOut351)>>1 ;
	end
end
FIFO  myfifo(.clk(clk) ,.reset(reset) ,.in(X) ,.out(oldData) ,.flag(flag));
medianFilterCell  m1(.X(X) ,.oldData(oldData) ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(0) ,.dataR_in(dataOut2) ,.dataL_in(0) 
	 ,.R_out(R1) ,.data_out(dataOut1)  );
medianFilterCell  m2(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R1) ,.dataR_in(dataOut3) ,.dataL_in(dataOut1) 
	 ,.R_out(R2) ,.data_out(dataOut2)  );
medianFilterCell  m3(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R2) ,.dataR_in(dataOut4) ,.dataL_in(dataOut2) 
	 ,.R_out(R3) ,.data_out(dataOut3)  );
medianFilterCell  m4(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R3) ,.dataR_in(dataOut5) ,.dataL_in(dataOut3) 
	 ,.R_out(R4) ,.data_out(dataOut4)  );
medianFilterCell  m5(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R4) ,.dataR_in(dataOut6) ,.dataL_in(dataOut4) 
	 ,.R_out(R5) ,.data_out(dataOut5)  );
medianFilterCell  m6(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R5) ,.dataR_in(dataOut7) ,.dataL_in(dataOut5) 
	 ,.R_out(R6) ,.data_out(dataOut6)  );
medianFilterCell  m7(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R6) ,.dataR_in(dataOut8) ,.dataL_in(dataOut6) 
	 ,.R_out(R7) ,.data_out(dataOut7)  );
medianFilterCell  m8(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R7) ,.dataR_in(dataOut9) ,.dataL_in(dataOut7) 
	 ,.R_out(R8) ,.data_out(dataOut8)  );
medianFilterCell  m9(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R8) ,.dataR_in(dataOut10) ,.dataL_in(dataOut8) 
	 ,.R_out(R9) ,.data_out(dataOut9)  );
medianFilterCell  m10(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R9) ,.dataR_in(dataOut11) ,.dataL_in(dataOut9) 
	 ,.R_out(R10) ,.data_out(dataOut10)  );
medianFilterCell  m11(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R10) ,.dataR_in(dataOut12) ,.dataL_in(dataOut10) 
	 ,.R_out(R11) ,.data_out(dataOut11)  );
medianFilterCell  m12(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R11) ,.dataR_in(dataOut13) ,.dataL_in(dataOut11) 
	 ,.R_out(R12) ,.data_out(dataOut12)  );
medianFilterCell  m13(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R12) ,.dataR_in(dataOut14) ,.dataL_in(dataOut12) 
	 ,.R_out(R13) ,.data_out(dataOut13)  );
medianFilterCell  m14(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R13) ,.dataR_in(dataOut15) ,.dataL_in(dataOut13) 
	 ,.R_out(R14) ,.data_out(dataOut14)  );
medianFilterCell  m15(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R14) ,.dataR_in(dataOut16) ,.dataL_in(dataOut14) 
	 ,.R_out(R15) ,.data_out(dataOut15)  );
medianFilterCell  m16(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R15) ,.dataR_in(dataOut17) ,.dataL_in(dataOut15) 
	 ,.R_out(R16) ,.data_out(dataOut16)  );
medianFilterCell  m17(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R16) ,.dataR_in(dataOut18) ,.dataL_in(dataOut16) 
	 ,.R_out(R17) ,.data_out(dataOut17)  );
medianFilterCell  m18(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R17) ,.dataR_in(dataOut19) ,.dataL_in(dataOut17) 
	 ,.R_out(R18) ,.data_out(dataOut18)  );
medianFilterCell  m19(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R18) ,.dataR_in(dataOut20) ,.dataL_in(dataOut18) 
	 ,.R_out(R19) ,.data_out(dataOut19)  );
medianFilterCell  m20(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R19) ,.dataR_in(dataOut21) ,.dataL_in(dataOut19) 
	 ,.R_out(R20) ,.data_out(dataOut20)  );
medianFilterCell  m21(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R20) ,.dataR_in(dataOut22) ,.dataL_in(dataOut20) 
	 ,.R_out(R21) ,.data_out(dataOut21)  );
medianFilterCell  m22(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R21) ,.dataR_in(dataOut23) ,.dataL_in(dataOut21) 
	 ,.R_out(R22) ,.data_out(dataOut22)  );
medianFilterCell  m23(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R22) ,.dataR_in(dataOut24) ,.dataL_in(dataOut22) 
	 ,.R_out(R23) ,.data_out(dataOut23)  );
medianFilterCell  m24(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R23) ,.dataR_in(dataOut25) ,.dataL_in(dataOut23) 
	 ,.R_out(R24) ,.data_out(dataOut24)  );
medianFilterCell  m25(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R24) ,.dataR_in(dataOut26) ,.dataL_in(dataOut24) 
	 ,.R_out(R25) ,.data_out(dataOut25)  );
medianFilterCell  m26(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R25) ,.dataR_in(dataOut27) ,.dataL_in(dataOut25) 
	 ,.R_out(R26) ,.data_out(dataOut26)  );
medianFilterCell  m27(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R26) ,.dataR_in(dataOut28) ,.dataL_in(dataOut26) 
	 ,.R_out(R27) ,.data_out(dataOut27)  );
medianFilterCell  m28(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R27) ,.dataR_in(dataOut29) ,.dataL_in(dataOut27) 
	 ,.R_out(R28) ,.data_out(dataOut28)  );
medianFilterCell  m29(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R28) ,.dataR_in(dataOut30) ,.dataL_in(dataOut28) 
	 ,.R_out(R29) ,.data_out(dataOut29)  );
medianFilterCell  m30(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R29) ,.dataR_in(dataOut31) ,.dataL_in(dataOut29) 
	 ,.R_out(R30) ,.data_out(dataOut30)  );
medianFilterCell  m31(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R30) ,.dataR_in(dataOut32) ,.dataL_in(dataOut30) 
	 ,.R_out(R31) ,.data_out(dataOut31)  );
medianFilterCell  m32(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R31) ,.dataR_in(dataOut33) ,.dataL_in(dataOut31) 
	 ,.R_out(R32) ,.data_out(dataOut32)  );
medianFilterCell  m33(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R32) ,.dataR_in(dataOut34) ,.dataL_in(dataOut32) 
	 ,.R_out(R33) ,.data_out(dataOut33)  );
medianFilterCell  m34(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R33) ,.dataR_in(dataOut35) ,.dataL_in(dataOut33) 
	 ,.R_out(R34) ,.data_out(dataOut34)  );
medianFilterCell  m35(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R34) ,.dataR_in(dataOut36) ,.dataL_in(dataOut34) 
	 ,.R_out(R35) ,.data_out(dataOut35)  );
medianFilterCell  m36(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R35) ,.dataR_in(dataOut37) ,.dataL_in(dataOut35) 
	 ,.R_out(R36) ,.data_out(dataOut36)  );
medianFilterCell  m37(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R36) ,.dataR_in(dataOut38) ,.dataL_in(dataOut36) 
	 ,.R_out(R37) ,.data_out(dataOut37)  );
medianFilterCell  m38(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R37) ,.dataR_in(dataOut39) ,.dataL_in(dataOut37) 
	 ,.R_out(R38) ,.data_out(dataOut38)  );
medianFilterCell  m39(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R38) ,.dataR_in(dataOut40) ,.dataL_in(dataOut38) 
	 ,.R_out(R39) ,.data_out(dataOut39)  );
medianFilterCell  m40(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R39) ,.dataR_in(dataOut41) ,.dataL_in(dataOut39) 
	 ,.R_out(R40) ,.data_out(dataOut40)  );
medianFilterCell  m41(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R40) ,.dataR_in(dataOut42) ,.dataL_in(dataOut40) 
	 ,.R_out(R41) ,.data_out(dataOut41)  );
medianFilterCell  m42(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R41) ,.dataR_in(dataOut43) ,.dataL_in(dataOut41) 
	 ,.R_out(R42) ,.data_out(dataOut42)  );
medianFilterCell  m43(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R42) ,.dataR_in(dataOut44) ,.dataL_in(dataOut42) 
	 ,.R_out(R43) ,.data_out(dataOut43)  );
medianFilterCell  m44(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R43) ,.dataR_in(dataOut45) ,.dataL_in(dataOut43) 
	 ,.R_out(R44) ,.data_out(dataOut44)  );
medianFilterCell  m45(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R44) ,.dataR_in(dataOut46) ,.dataL_in(dataOut44) 
	 ,.R_out(R45) ,.data_out(dataOut45)  );
medianFilterCell  m46(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R45) ,.dataR_in(dataOut47) ,.dataL_in(dataOut45) 
	 ,.R_out(R46) ,.data_out(dataOut46)  );
medianFilterCell  m47(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R46) ,.dataR_in(dataOut48) ,.dataL_in(dataOut46) 
	 ,.R_out(R47) ,.data_out(dataOut47)  );
medianFilterCell  m48(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R47) ,.dataR_in(dataOut49) ,.dataL_in(dataOut47) 
	 ,.R_out(R48) ,.data_out(dataOut48)  );
medianFilterCell  m49(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R48) ,.dataR_in(dataOut50) ,.dataL_in(dataOut48) 
	 ,.R_out(R49) ,.data_out(dataOut49)  );
medianFilterCell  m50(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R49) ,.dataR_in(dataOut51) ,.dataL_in(dataOut49) 
	 ,.R_out(R50) ,.data_out(dataOut50)  );
medianFilterCell  m51(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R50) ,.dataR_in(dataOut52) ,.dataL_in(dataOut50) 
	 ,.R_out(R51) ,.data_out(dataOut51)  );
medianFilterCell  m52(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R51) ,.dataR_in(dataOut53) ,.dataL_in(dataOut51) 
	 ,.R_out(R52) ,.data_out(dataOut52)  );
medianFilterCell  m53(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R52) ,.dataR_in(dataOut54) ,.dataL_in(dataOut52) 
	 ,.R_out(R53) ,.data_out(dataOut53)  );
medianFilterCell  m54(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R53) ,.dataR_in(dataOut55) ,.dataL_in(dataOut53) 
	 ,.R_out(R54) ,.data_out(dataOut54)  );
medianFilterCell  m55(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R54) ,.dataR_in(dataOut56) ,.dataL_in(dataOut54) 
	 ,.R_out(R55) ,.data_out(dataOut55)  );
medianFilterCell  m56(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R55) ,.dataR_in(dataOut57) ,.dataL_in(dataOut55) 
	 ,.R_out(R56) ,.data_out(dataOut56)  );
medianFilterCell  m57(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R56) ,.dataR_in(dataOut58) ,.dataL_in(dataOut56) 
	 ,.R_out(R57) ,.data_out(dataOut57)  );
medianFilterCell  m58(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R57) ,.dataR_in(dataOut59) ,.dataL_in(dataOut57) 
	 ,.R_out(R58) ,.data_out(dataOut58)  );
medianFilterCell  m59(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R58) ,.dataR_in(dataOut60) ,.dataL_in(dataOut58) 
	 ,.R_out(R59) ,.data_out(dataOut59)  );
medianFilterCell  m60(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R59) ,.dataR_in(dataOut61) ,.dataL_in(dataOut59) 
	 ,.R_out(R60) ,.data_out(dataOut60)  );
medianFilterCell  m61(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R60) ,.dataR_in(dataOut62) ,.dataL_in(dataOut60) 
	 ,.R_out(R61) ,.data_out(dataOut61)  );
medianFilterCell  m62(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R61) ,.dataR_in(dataOut63) ,.dataL_in(dataOut61) 
	 ,.R_out(R62) ,.data_out(dataOut62)  );
medianFilterCell  m63(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R62) ,.dataR_in(dataOut64) ,.dataL_in(dataOut62) 
	 ,.R_out(R63) ,.data_out(dataOut63)  );
medianFilterCell  m64(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R63) ,.dataR_in(dataOut65) ,.dataL_in(dataOut63) 
	 ,.R_out(R64) ,.data_out(dataOut64)  );
medianFilterCell  m65(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R64) ,.dataR_in(dataOut66) ,.dataL_in(dataOut64) 
	 ,.R_out(R65) ,.data_out(dataOut65)  );
medianFilterCell  m66(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R65) ,.dataR_in(dataOut67) ,.dataL_in(dataOut65) 
	 ,.R_out(R66) ,.data_out(dataOut66)  );
medianFilterCell  m67(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R66) ,.dataR_in(dataOut68) ,.dataL_in(dataOut66) 
	 ,.R_out(R67) ,.data_out(dataOut67)  );
medianFilterCell  m68(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R67) ,.dataR_in(dataOut69) ,.dataL_in(dataOut67) 
	 ,.R_out(R68) ,.data_out(dataOut68)  );
medianFilterCell  m69(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R68) ,.dataR_in(dataOut70) ,.dataL_in(dataOut68) 
	 ,.R_out(R69) ,.data_out(dataOut69)  );
medianFilterCell  m70(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R69) ,.dataR_in(dataOut71) ,.dataL_in(dataOut69) 
	 ,.R_out(R70) ,.data_out(dataOut70)  );
medianFilterCell  m71(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R70) ,.dataR_in(dataOut72) ,.dataL_in(dataOut70) 
	 ,.R_out(R71) ,.data_out(dataOut71)  );
medianFilterCell  m72(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R71) ,.dataR_in(dataOut73) ,.dataL_in(dataOut71) 
	 ,.R_out(R72) ,.data_out(dataOut72)  );
medianFilterCell  m73(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R72) ,.dataR_in(dataOut74) ,.dataL_in(dataOut72) 
	 ,.R_out(R73) ,.data_out(dataOut73)  );
medianFilterCell  m74(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R73) ,.dataR_in(dataOut75) ,.dataL_in(dataOut73) 
	 ,.R_out(R74) ,.data_out(dataOut74)  );
medianFilterCell  m75(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R74) ,.dataR_in(dataOut76) ,.dataL_in(dataOut74) 
	 ,.R_out(R75) ,.data_out(dataOut75)  );
medianFilterCell  m76(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R75) ,.dataR_in(dataOut77) ,.dataL_in(dataOut75) 
	 ,.R_out(R76) ,.data_out(dataOut76)  );
medianFilterCell  m77(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R76) ,.dataR_in(dataOut78) ,.dataL_in(dataOut76) 
	 ,.R_out(R77) ,.data_out(dataOut77)  );
medianFilterCell  m78(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R77) ,.dataR_in(dataOut79) ,.dataL_in(dataOut77) 
	 ,.R_out(R78) ,.data_out(dataOut78)  );
medianFilterCell  m79(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R78) ,.dataR_in(dataOut80) ,.dataL_in(dataOut78) 
	 ,.R_out(R79) ,.data_out(dataOut79)  );
medianFilterCell  m80(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R79) ,.dataR_in(dataOut81) ,.dataL_in(dataOut79) 
	 ,.R_out(R80) ,.data_out(dataOut80)  );
medianFilterCell  m81(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R80) ,.dataR_in(dataOut82) ,.dataL_in(dataOut80) 
	 ,.R_out(R81) ,.data_out(dataOut81)  );
medianFilterCell  m82(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R81) ,.dataR_in(dataOut83) ,.dataL_in(dataOut81) 
	 ,.R_out(R82) ,.data_out(dataOut82)  );
medianFilterCell  m83(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R82) ,.dataR_in(dataOut84) ,.dataL_in(dataOut82) 
	 ,.R_out(R83) ,.data_out(dataOut83)  );
medianFilterCell  m84(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R83) ,.dataR_in(dataOut85) ,.dataL_in(dataOut83) 
	 ,.R_out(R84) ,.data_out(dataOut84)  );
medianFilterCell  m85(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R84) ,.dataR_in(dataOut86) ,.dataL_in(dataOut84) 
	 ,.R_out(R85) ,.data_out(dataOut85)  );
medianFilterCell  m86(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R85) ,.dataR_in(dataOut87) ,.dataL_in(dataOut85) 
	 ,.R_out(R86) ,.data_out(dataOut86)  );
medianFilterCell  m87(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R86) ,.dataR_in(dataOut88) ,.dataL_in(dataOut86) 
	 ,.R_out(R87) ,.data_out(dataOut87)  );
medianFilterCell  m88(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R87) ,.dataR_in(dataOut89) ,.dataL_in(dataOut87) 
	 ,.R_out(R88) ,.data_out(dataOut88)  );
medianFilterCell  m89(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R88) ,.dataR_in(dataOut90) ,.dataL_in(dataOut88) 
	 ,.R_out(R89) ,.data_out(dataOut89)  );
medianFilterCell  m90(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R89) ,.dataR_in(dataOut91) ,.dataL_in(dataOut89) 
	 ,.R_out(R90) ,.data_out(dataOut90)  );
medianFilterCell  m91(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R90) ,.dataR_in(dataOut92) ,.dataL_in(dataOut90) 
	 ,.R_out(R91) ,.data_out(dataOut91)  );
medianFilterCell  m92(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R91) ,.dataR_in(dataOut93) ,.dataL_in(dataOut91) 
	 ,.R_out(R92) ,.data_out(dataOut92)  );
medianFilterCell  m93(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R92) ,.dataR_in(dataOut94) ,.dataL_in(dataOut92) 
	 ,.R_out(R93) ,.data_out(dataOut93)  );
medianFilterCell  m94(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R93) ,.dataR_in(dataOut95) ,.dataL_in(dataOut93) 
	 ,.R_out(R94) ,.data_out(dataOut94)  );
medianFilterCell  m95(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R94) ,.dataR_in(dataOut96) ,.dataL_in(dataOut94) 
	 ,.R_out(R95) ,.data_out(dataOut95)  );
medianFilterCell  m96(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R95) ,.dataR_in(dataOut97) ,.dataL_in(dataOut95) 
	 ,.R_out(R96) ,.data_out(dataOut96)  );
medianFilterCell  m97(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R96) ,.dataR_in(dataOut98) ,.dataL_in(dataOut96) 
	 ,.R_out(R97) ,.data_out(dataOut97)  );
medianFilterCell  m98(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R97) ,.dataR_in(dataOut99) ,.dataL_in(dataOut97) 
	 ,.R_out(R98) ,.data_out(dataOut98)  );
medianFilterCell  m99(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R98) ,.dataR_in(dataOut100) ,.dataL_in(dataOut98) 
	 ,.R_out(R99) ,.data_out(dataOut99)  );
medianFilterCell  m100(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R99) ,.dataR_in(dataOut101) ,.dataL_in(dataOut99) 
	 ,.R_out(R100) ,.data_out(dataOut100)  );
medianFilterCell  m101(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R100) ,.dataR_in(dataOut102) ,.dataL_in(dataOut100) 
	 ,.R_out(R101) ,.data_out(dataOut101)  );
medianFilterCell  m102(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R101) ,.dataR_in(dataOut103) ,.dataL_in(dataOut101) 
	 ,.R_out(R102) ,.data_out(dataOut102)  );
medianFilterCell  m103(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R102) ,.dataR_in(dataOut104) ,.dataL_in(dataOut102) 
	 ,.R_out(R103) ,.data_out(dataOut103)  );
medianFilterCell  m104(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R103) ,.dataR_in(dataOut105) ,.dataL_in(dataOut103) 
	 ,.R_out(R104) ,.data_out(dataOut104)  );
medianFilterCell  m105(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R104) ,.dataR_in(dataOut106) ,.dataL_in(dataOut104) 
	 ,.R_out(R105) ,.data_out(dataOut105)  );
medianFilterCell  m106(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R105) ,.dataR_in(dataOut107) ,.dataL_in(dataOut105) 
	 ,.R_out(R106) ,.data_out(dataOut106)  );
medianFilterCell  m107(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R106) ,.dataR_in(dataOut108) ,.dataL_in(dataOut106) 
	 ,.R_out(R107) ,.data_out(dataOut107)  );
medianFilterCell  m108(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R107) ,.dataR_in(dataOut109) ,.dataL_in(dataOut107) 
	 ,.R_out(R108) ,.data_out(dataOut108)  );
medianFilterCell  m109(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R108) ,.dataR_in(dataOut110) ,.dataL_in(dataOut108) 
	 ,.R_out(R109) ,.data_out(dataOut109)  );
medianFilterCell  m110(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R109) ,.dataR_in(dataOut111) ,.dataL_in(dataOut109) 
	 ,.R_out(R110) ,.data_out(dataOut110)  );
medianFilterCell  m111(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R110) ,.dataR_in(dataOut112) ,.dataL_in(dataOut110) 
	 ,.R_out(R111) ,.data_out(dataOut111)  );
medianFilterCell  m112(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R111) ,.dataR_in(dataOut113) ,.dataL_in(dataOut111) 
	 ,.R_out(R112) ,.data_out(dataOut112)  );
medianFilterCell  m113(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R112) ,.dataR_in(dataOut114) ,.dataL_in(dataOut112) 
	 ,.R_out(R113) ,.data_out(dataOut113)  );
medianFilterCell  m114(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R113) ,.dataR_in(dataOut115) ,.dataL_in(dataOut113) 
	 ,.R_out(R114) ,.data_out(dataOut114)  );
medianFilterCell  m115(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R114) ,.dataR_in(dataOut116) ,.dataL_in(dataOut114) 
	 ,.R_out(R115) ,.data_out(dataOut115)  );
medianFilterCell  m116(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R115) ,.dataR_in(dataOut117) ,.dataL_in(dataOut115) 
	 ,.R_out(R116) ,.data_out(dataOut116)  );
medianFilterCell  m117(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R116) ,.dataR_in(dataOut118) ,.dataL_in(dataOut116) 
	 ,.R_out(R117) ,.data_out(dataOut117)  );
medianFilterCell  m118(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R117) ,.dataR_in(dataOut119) ,.dataL_in(dataOut117) 
	 ,.R_out(R118) ,.data_out(dataOut118)  );
medianFilterCell  m119(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R118) ,.dataR_in(dataOut120) ,.dataL_in(dataOut118) 
	 ,.R_out(R119) ,.data_out(dataOut119)  );
medianFilterCell  m120(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R119) ,.dataR_in(dataOut121) ,.dataL_in(dataOut119) 
	 ,.R_out(R120) ,.data_out(dataOut120)  );
medianFilterCell  m121(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R120) ,.dataR_in(dataOut122) ,.dataL_in(dataOut120) 
	 ,.R_out(R121) ,.data_out(dataOut121)  );
medianFilterCell  m122(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R121) ,.dataR_in(dataOut123) ,.dataL_in(dataOut121) 
	 ,.R_out(R122) ,.data_out(dataOut122)  );
medianFilterCell  m123(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R122) ,.dataR_in(dataOut124) ,.dataL_in(dataOut122) 
	 ,.R_out(R123) ,.data_out(dataOut123)  );
medianFilterCell  m124(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R123) ,.dataR_in(dataOut125) ,.dataL_in(dataOut123) 
	 ,.R_out(R124) ,.data_out(dataOut124)  );
medianFilterCell  m125(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R124) ,.dataR_in(dataOut126) ,.dataL_in(dataOut124) 
	 ,.R_out(R125) ,.data_out(dataOut125)  );
medianFilterCell  m126(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R125) ,.dataR_in(dataOut127) ,.dataL_in(dataOut125) 
	 ,.R_out(R126) ,.data_out(dataOut126)  );
medianFilterCell  m127(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R126) ,.dataR_in(dataOut128) ,.dataL_in(dataOut126) 
	 ,.R_out(R127) ,.data_out(dataOut127)  );
medianFilterCell  m128(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R127) ,.dataR_in(dataOut129) ,.dataL_in(dataOut127) 
	 ,.R_out(R128) ,.data_out(dataOut128)  );
medianFilterCell  m129(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R128) ,.dataR_in(dataOut130) ,.dataL_in(dataOut128) 
	 ,.R_out(R129) ,.data_out(dataOut129)  );
medianFilterCell  m130(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R129) ,.dataR_in(dataOut131) ,.dataL_in(dataOut129) 
	 ,.R_out(R130) ,.data_out(dataOut130)  );
medianFilterCell  m131(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R130) ,.dataR_in(dataOut132) ,.dataL_in(dataOut130) 
	 ,.R_out(R131) ,.data_out(dataOut131)  );
medianFilterCell  m132(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R131) ,.dataR_in(dataOut133) ,.dataL_in(dataOut131) 
	 ,.R_out(R132) ,.data_out(dataOut132)  );
medianFilterCell  m133(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R132) ,.dataR_in(dataOut134) ,.dataL_in(dataOut132) 
	 ,.R_out(R133) ,.data_out(dataOut133)  );
medianFilterCell  m134(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R133) ,.dataR_in(dataOut135) ,.dataL_in(dataOut133) 
	 ,.R_out(R134) ,.data_out(dataOut134)  );
medianFilterCell  m135(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R134) ,.dataR_in(dataOut136) ,.dataL_in(dataOut134) 
	 ,.R_out(R135) ,.data_out(dataOut135)  );
medianFilterCell  m136(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R135) ,.dataR_in(dataOut137) ,.dataL_in(dataOut135) 
	 ,.R_out(R136) ,.data_out(dataOut136)  );
medianFilterCell  m137(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R136) ,.dataR_in(dataOut138) ,.dataL_in(dataOut136) 
	 ,.R_out(R137) ,.data_out(dataOut137)  );
medianFilterCell  m138(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R137) ,.dataR_in(dataOut139) ,.dataL_in(dataOut137) 
	 ,.R_out(R138) ,.data_out(dataOut138)  );
medianFilterCell  m139(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R138) ,.dataR_in(dataOut140) ,.dataL_in(dataOut138) 
	 ,.R_out(R139) ,.data_out(dataOut139)  );
medianFilterCell  m140(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R139) ,.dataR_in(dataOut141) ,.dataL_in(dataOut139) 
	 ,.R_out(R140) ,.data_out(dataOut140)  );
medianFilterCell  m141(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R140) ,.dataR_in(dataOut142) ,.dataL_in(dataOut140) 
	 ,.R_out(R141) ,.data_out(dataOut141)  );
medianFilterCell  m142(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R141) ,.dataR_in(dataOut143) ,.dataL_in(dataOut141) 
	 ,.R_out(R142) ,.data_out(dataOut142)  );
medianFilterCell  m143(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R142) ,.dataR_in(dataOut144) ,.dataL_in(dataOut142) 
	 ,.R_out(R143) ,.data_out(dataOut143)  );
medianFilterCell  m144(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R143) ,.dataR_in(dataOut145) ,.dataL_in(dataOut143) 
	 ,.R_out(R144) ,.data_out(dataOut144)  );
medianFilterCell  m145(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R144) ,.dataR_in(dataOut146) ,.dataL_in(dataOut144) 
	 ,.R_out(R145) ,.data_out(dataOut145)  );
medianFilterCell  m146(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R145) ,.dataR_in(dataOut147) ,.dataL_in(dataOut145) 
	 ,.R_out(R146) ,.data_out(dataOut146)  );
medianFilterCell  m147(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R146) ,.dataR_in(dataOut148) ,.dataL_in(dataOut146) 
	 ,.R_out(R147) ,.data_out(dataOut147)  );
medianFilterCell  m148(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R147) ,.dataR_in(dataOut149) ,.dataL_in(dataOut147) 
	 ,.R_out(R148) ,.data_out(dataOut148)  );
medianFilterCell  m149(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R148) ,.dataR_in(dataOut150) ,.dataL_in(dataOut148) 
	 ,.R_out(R149) ,.data_out(dataOut149)  );
medianFilterCell  m150(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R149) ,.dataR_in(dataOut151) ,.dataL_in(dataOut149) 
	 ,.R_out(R150) ,.data_out(dataOut150)  );
medianFilterCell  m151(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R150) ,.dataR_in(dataOut152) ,.dataL_in(dataOut150) 
	 ,.R_out(R151) ,.data_out(dataOut151)  );
medianFilterCell  m152(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R151) ,.dataR_in(dataOut153) ,.dataL_in(dataOut151) 
	 ,.R_out(R152) ,.data_out(dataOut152)  );
medianFilterCell  m153(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R152) ,.dataR_in(dataOut154) ,.dataL_in(dataOut152) 
	 ,.R_out(R153) ,.data_out(dataOut153)  );
medianFilterCell  m154(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R153) ,.dataR_in(dataOut155) ,.dataL_in(dataOut153) 
	 ,.R_out(R154) ,.data_out(dataOut154)  );
medianFilterCell  m155(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R154) ,.dataR_in(dataOut156) ,.dataL_in(dataOut154) 
	 ,.R_out(R155) ,.data_out(dataOut155)  );
medianFilterCell  m156(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R155) ,.dataR_in(dataOut157) ,.dataL_in(dataOut155) 
	 ,.R_out(R156) ,.data_out(dataOut156)  );
medianFilterCell  m157(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R156) ,.dataR_in(dataOut158) ,.dataL_in(dataOut156) 
	 ,.R_out(R157) ,.data_out(dataOut157)  );
medianFilterCell  m158(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R157) ,.dataR_in(dataOut159) ,.dataL_in(dataOut157) 
	 ,.R_out(R158) ,.data_out(dataOut158)  );
medianFilterCell  m159(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R158) ,.dataR_in(dataOut160) ,.dataL_in(dataOut158) 
	 ,.R_out(R159) ,.data_out(dataOut159)  );
medianFilterCell  m160(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R159) ,.dataR_in(dataOut161) ,.dataL_in(dataOut159) 
	 ,.R_out(R160) ,.data_out(dataOut160)  );
medianFilterCell  m161(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R160) ,.dataR_in(dataOut162) ,.dataL_in(dataOut160) 
	 ,.R_out(R161) ,.data_out(dataOut161)  );
medianFilterCell  m162(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R161) ,.dataR_in(dataOut163) ,.dataL_in(dataOut161) 
	 ,.R_out(R162) ,.data_out(dataOut162)  );
medianFilterCell  m163(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R162) ,.dataR_in(dataOut164) ,.dataL_in(dataOut162) 
	 ,.R_out(R163) ,.data_out(dataOut163)  );
medianFilterCell  m164(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R163) ,.dataR_in(dataOut165) ,.dataL_in(dataOut163) 
	 ,.R_out(R164) ,.data_out(dataOut164)  );
medianFilterCell  m165(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R164) ,.dataR_in(dataOut166) ,.dataL_in(dataOut164) 
	 ,.R_out(R165) ,.data_out(dataOut165)  );
medianFilterCell  m166(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R165) ,.dataR_in(dataOut167) ,.dataL_in(dataOut165) 
	 ,.R_out(R166) ,.data_out(dataOut166)  );
medianFilterCell  m167(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R166) ,.dataR_in(dataOut168) ,.dataL_in(dataOut166) 
	 ,.R_out(R167) ,.data_out(dataOut167)  );
medianFilterCell  m168(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R167) ,.dataR_in(dataOut169) ,.dataL_in(dataOut167) 
	 ,.R_out(R168) ,.data_out(dataOut168)  );
medianFilterCell  m169(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R168) ,.dataR_in(dataOut170) ,.dataL_in(dataOut168) 
	 ,.R_out(R169) ,.data_out(dataOut169)  );
medianFilterCell  m170(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R169) ,.dataR_in(dataOut171) ,.dataL_in(dataOut169) 
	 ,.R_out(R170) ,.data_out(dataOut170)  );
medianFilterCell  m171(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R170) ,.dataR_in(dataOut172) ,.dataL_in(dataOut170) 
	 ,.R_out(R171) ,.data_out(dataOut171)  );
medianFilterCell  m172(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R171) ,.dataR_in(dataOut173) ,.dataL_in(dataOut171) 
	 ,.R_out(R172) ,.data_out(dataOut172)  );
medianFilterCell  m173(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R172) ,.dataR_in(dataOut174) ,.dataL_in(dataOut172) 
	 ,.R_out(R173) ,.data_out(dataOut173)  );
medianFilterCell  m174(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R173) ,.dataR_in(dataOut175) ,.dataL_in(dataOut173) 
	 ,.R_out(R174) ,.data_out(dataOut174)  );
medianFilterCell  m175(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R174) ,.dataR_in(dataOut176) ,.dataL_in(dataOut174) 
	 ,.R_out(R175) ,.data_out(dataOut175)  );
medianFilterCell  m176(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R175) ,.dataR_in(dataOut177) ,.dataL_in(dataOut175) 
	 ,.R_out(R176) ,.data_out(dataOut176)  );
medianFilterCell  m177(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R176) ,.dataR_in(dataOut178) ,.dataL_in(dataOut176) 
	 ,.R_out(R177) ,.data_out(dataOut177)  );
medianFilterCell  m178(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R177) ,.dataR_in(dataOut179) ,.dataL_in(dataOut177) 
	 ,.R_out(R178) ,.data_out(dataOut178)  );
medianFilterCell  m179(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R178) ,.dataR_in(dataOut180) ,.dataL_in(dataOut178) 
	 ,.R_out(R179) ,.data_out(dataOut179)  );
medianFilterCell  m180(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R179) ,.dataR_in(dataOut181) ,.dataL_in(dataOut179) 
	 ,.R_out(R180) ,.data_out(dataOut180)  );
medianFilterCell  m181(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R180) ,.dataR_in(dataOut182) ,.dataL_in(dataOut180) 
	 ,.R_out(R181) ,.data_out(dataOut181)  );
medianFilterCell  m182(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R181) ,.dataR_in(dataOut183) ,.dataL_in(dataOut181) 
	 ,.R_out(R182) ,.data_out(dataOut182)  );
medianFilterCell  m183(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R182) ,.dataR_in(dataOut184) ,.dataL_in(dataOut182) 
	 ,.R_out(R183) ,.data_out(dataOut183)  );
medianFilterCell  m184(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R183) ,.dataR_in(dataOut185) ,.dataL_in(dataOut183) 
	 ,.R_out(R184) ,.data_out(dataOut184)  );
medianFilterCell  m185(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R184) ,.dataR_in(dataOut186) ,.dataL_in(dataOut184) 
	 ,.R_out(R185) ,.data_out(dataOut185)  );
medianFilterCell  m186(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R185) ,.dataR_in(dataOut187) ,.dataL_in(dataOut185) 
	 ,.R_out(R186) ,.data_out(dataOut186)  );
medianFilterCell  m187(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R186) ,.dataR_in(dataOut188) ,.dataL_in(dataOut186) 
	 ,.R_out(R187) ,.data_out(dataOut187)  );
medianFilterCell  m188(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R187) ,.dataR_in(dataOut189) ,.dataL_in(dataOut187) 
	 ,.R_out(R188) ,.data_out(dataOut188)  );
medianFilterCell  m189(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R188) ,.dataR_in(dataOut190) ,.dataL_in(dataOut188) 
	 ,.R_out(R189) ,.data_out(dataOut189)  );
medianFilterCell  m190(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R189) ,.dataR_in(dataOut191) ,.dataL_in(dataOut189) 
	 ,.R_out(R190) ,.data_out(dataOut190)  );
medianFilterCell  m191(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R190) ,.dataR_in(dataOut192) ,.dataL_in(dataOut190) 
	 ,.R_out(R191) ,.data_out(dataOut191)  );
medianFilterCell  m192(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R191) ,.dataR_in(dataOut193) ,.dataL_in(dataOut191) 
	 ,.R_out(R192) ,.data_out(dataOut192)  );
medianFilterCell  m193(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R192) ,.dataR_in(dataOut194) ,.dataL_in(dataOut192) 
	 ,.R_out(R193) ,.data_out(dataOut193)  );
medianFilterCell  m194(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R193) ,.dataR_in(dataOut195) ,.dataL_in(dataOut193) 
	 ,.R_out(R194) ,.data_out(dataOut194)  );
medianFilterCell  m195(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R194) ,.dataR_in(dataOut196) ,.dataL_in(dataOut194) 
	 ,.R_out(R195) ,.data_out(dataOut195)  );
medianFilterCell  m196(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R195) ,.dataR_in(dataOut197) ,.dataL_in(dataOut195) 
	 ,.R_out(R196) ,.data_out(dataOut196)  );
medianFilterCell  m197(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R196) ,.dataR_in(dataOut198) ,.dataL_in(dataOut196) 
	 ,.R_out(R197) ,.data_out(dataOut197)  );
medianFilterCell  m198(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R197) ,.dataR_in(dataOut199) ,.dataL_in(dataOut197) 
	 ,.R_out(R198) ,.data_out(dataOut198)  );
medianFilterCell  m199(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R198) ,.dataR_in(dataOut200) ,.dataL_in(dataOut198) 
	 ,.R_out(R199) ,.data_out(dataOut199)  );
medianFilterCell  m200(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R199) ,.dataR_in(dataOut201) ,.dataL_in(dataOut199) 
	 ,.R_out(R200) ,.data_out(dataOut200)  );
medianFilterCell  m201(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R200) ,.dataR_in(dataOut202) ,.dataL_in(dataOut200) 
	 ,.R_out(R201) ,.data_out(dataOut201)  );
medianFilterCell  m202(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R201) ,.dataR_in(dataOut203) ,.dataL_in(dataOut201) 
	 ,.R_out(R202) ,.data_out(dataOut202)  );
medianFilterCell  m203(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R202) ,.dataR_in(dataOut204) ,.dataL_in(dataOut202) 
	 ,.R_out(R203) ,.data_out(dataOut203)  );
medianFilterCell  m204(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R203) ,.dataR_in(dataOut205) ,.dataL_in(dataOut203) 
	 ,.R_out(R204) ,.data_out(dataOut204)  );
medianFilterCell  m205(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R204) ,.dataR_in(dataOut206) ,.dataL_in(dataOut204) 
	 ,.R_out(R205) ,.data_out(dataOut205)  );
medianFilterCell  m206(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R205) ,.dataR_in(dataOut207) ,.dataL_in(dataOut205) 
	 ,.R_out(R206) ,.data_out(dataOut206)  );
medianFilterCell  m207(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R206) ,.dataR_in(dataOut208) ,.dataL_in(dataOut206) 
	 ,.R_out(R207) ,.data_out(dataOut207)  );
medianFilterCell  m208(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R207) ,.dataR_in(dataOut209) ,.dataL_in(dataOut207) 
	 ,.R_out(R208) ,.data_out(dataOut208)  );
medianFilterCell  m209(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R208) ,.dataR_in(dataOut210) ,.dataL_in(dataOut208) 
	 ,.R_out(R209) ,.data_out(dataOut209)  );
medianFilterCell  m210(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R209) ,.dataR_in(dataOut211) ,.dataL_in(dataOut209) 
	 ,.R_out(R210) ,.data_out(dataOut210)  );
medianFilterCell  m211(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R210) ,.dataR_in(dataOut212) ,.dataL_in(dataOut210) 
	 ,.R_out(R211) ,.data_out(dataOut211)  );
medianFilterCell  m212(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R211) ,.dataR_in(dataOut213) ,.dataL_in(dataOut211) 
	 ,.R_out(R212) ,.data_out(dataOut212)  );
medianFilterCell  m213(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R212) ,.dataR_in(dataOut214) ,.dataL_in(dataOut212) 
	 ,.R_out(R213) ,.data_out(dataOut213)  );
medianFilterCell  m214(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R213) ,.dataR_in(dataOut215) ,.dataL_in(dataOut213) 
	 ,.R_out(R214) ,.data_out(dataOut214)  );
medianFilterCell  m215(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R214) ,.dataR_in(dataOut216) ,.dataL_in(dataOut214) 
	 ,.R_out(R215) ,.data_out(dataOut215)  );
medianFilterCell  m216(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R215) ,.dataR_in(dataOut217) ,.dataL_in(dataOut215) 
	 ,.R_out(R216) ,.data_out(dataOut216)  );
medianFilterCell  m217(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R216) ,.dataR_in(dataOut218) ,.dataL_in(dataOut216) 
	 ,.R_out(R217) ,.data_out(dataOut217)  );
medianFilterCell  m218(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R217) ,.dataR_in(dataOut219) ,.dataL_in(dataOut217) 
	 ,.R_out(R218) ,.data_out(dataOut218)  );
medianFilterCell  m219(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R218) ,.dataR_in(dataOut220) ,.dataL_in(dataOut218) 
	 ,.R_out(R219) ,.data_out(dataOut219)  );
medianFilterCell  m220(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R219) ,.dataR_in(dataOut221) ,.dataL_in(dataOut219) 
	 ,.R_out(R220) ,.data_out(dataOut220)  );
medianFilterCell  m221(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R220) ,.dataR_in(dataOut222) ,.dataL_in(dataOut220) 
	 ,.R_out(R221) ,.data_out(dataOut221)  );
medianFilterCell  m222(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R221) ,.dataR_in(dataOut223) ,.dataL_in(dataOut221) 
	 ,.R_out(R222) ,.data_out(dataOut222)  );
medianFilterCell  m223(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R222) ,.dataR_in(dataOut224) ,.dataL_in(dataOut222) 
	 ,.R_out(R223) ,.data_out(dataOut223)  );
medianFilterCell  m224(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R223) ,.dataR_in(dataOut225) ,.dataL_in(dataOut223) 
	 ,.R_out(R224) ,.data_out(dataOut224)  );
medianFilterCell  m225(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R224) ,.dataR_in(dataOut226) ,.dataL_in(dataOut224) 
	 ,.R_out(R225) ,.data_out(dataOut225)  );
medianFilterCell  m226(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R225) ,.dataR_in(dataOut227) ,.dataL_in(dataOut225) 
	 ,.R_out(R226) ,.data_out(dataOut226)  );
medianFilterCell  m227(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R226) ,.dataR_in(dataOut228) ,.dataL_in(dataOut226) 
	 ,.R_out(R227) ,.data_out(dataOut227)  );
medianFilterCell  m228(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R227) ,.dataR_in(dataOut229) ,.dataL_in(dataOut227) 
	 ,.R_out(R228) ,.data_out(dataOut228)  );
medianFilterCell  m229(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R228) ,.dataR_in(dataOut230) ,.dataL_in(dataOut228) 
	 ,.R_out(R229) ,.data_out(dataOut229)  );
medianFilterCell  m230(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R229) ,.dataR_in(dataOut231) ,.dataL_in(dataOut229) 
	 ,.R_out(R230) ,.data_out(dataOut230)  );
medianFilterCell  m231(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R230) ,.dataR_in(dataOut232) ,.dataL_in(dataOut230) 
	 ,.R_out(R231) ,.data_out(dataOut231)  );
medianFilterCell  m232(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R231) ,.dataR_in(dataOut233) ,.dataL_in(dataOut231) 
	 ,.R_out(R232) ,.data_out(dataOut232)  );
medianFilterCell  m233(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R232) ,.dataR_in(dataOut234) ,.dataL_in(dataOut232) 
	 ,.R_out(R233) ,.data_out(dataOut233)  );
medianFilterCell  m234(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R233) ,.dataR_in(dataOut235) ,.dataL_in(dataOut233) 
	 ,.R_out(R234) ,.data_out(dataOut234)  );
medianFilterCell  m235(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R234) ,.dataR_in(dataOut236) ,.dataL_in(dataOut234) 
	 ,.R_out(R235) ,.data_out(dataOut235)  );
medianFilterCell  m236(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R235) ,.dataR_in(dataOut237) ,.dataL_in(dataOut235) 
	 ,.R_out(R236) ,.data_out(dataOut236)  );
medianFilterCell  m237(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R236) ,.dataR_in(dataOut238) ,.dataL_in(dataOut236) 
	 ,.R_out(R237) ,.data_out(dataOut237)  );
medianFilterCell  m238(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R237) ,.dataR_in(dataOut239) ,.dataL_in(dataOut237) 
	 ,.R_out(R238) ,.data_out(dataOut238)  );
medianFilterCell  m239(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R238) ,.dataR_in(dataOut240) ,.dataL_in(dataOut238) 
	 ,.R_out(R239) ,.data_out(dataOut239)  );
medianFilterCell  m240(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R239) ,.dataR_in(dataOut241) ,.dataL_in(dataOut239) 
	 ,.R_out(R240) ,.data_out(dataOut240)  );
medianFilterCell  m241(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R240) ,.dataR_in(dataOut242) ,.dataL_in(dataOut240) 
	 ,.R_out(R241) ,.data_out(dataOut241)  );
medianFilterCell  m242(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R241) ,.dataR_in(dataOut243) ,.dataL_in(dataOut241) 
	 ,.R_out(R242) ,.data_out(dataOut242)  );
medianFilterCell  m243(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R242) ,.dataR_in(dataOut244) ,.dataL_in(dataOut242) 
	 ,.R_out(R243) ,.data_out(dataOut243)  );
medianFilterCell  m244(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R243) ,.dataR_in(dataOut245) ,.dataL_in(dataOut243) 
	 ,.R_out(R244) ,.data_out(dataOut244)  );
medianFilterCell  m245(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R244) ,.dataR_in(dataOut246) ,.dataL_in(dataOut244) 
	 ,.R_out(R245) ,.data_out(dataOut245)  );
medianFilterCell  m246(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R245) ,.dataR_in(dataOut247) ,.dataL_in(dataOut245) 
	 ,.R_out(R246) ,.data_out(dataOut246)  );
medianFilterCell  m247(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R246) ,.dataR_in(dataOut248) ,.dataL_in(dataOut246) 
	 ,.R_out(R247) ,.data_out(dataOut247)  );
medianFilterCell  m248(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R247) ,.dataR_in(dataOut249) ,.dataL_in(dataOut247) 
	 ,.R_out(R248) ,.data_out(dataOut248)  );
medianFilterCell  m249(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R248) ,.dataR_in(dataOut250) ,.dataL_in(dataOut248) 
	 ,.R_out(R249) ,.data_out(dataOut249)  );
medianFilterCell  m250(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R249) ,.dataR_in(dataOut251) ,.dataL_in(dataOut249) 
	 ,.R_out(R250) ,.data_out(dataOut250)  );
medianFilterCell  m251(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R250) ,.dataR_in(dataOut252) ,.dataL_in(dataOut250) 
	 ,.R_out(R251) ,.data_out(dataOut251)  );
medianFilterCell  m252(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R251) ,.dataR_in(dataOut253) ,.dataL_in(dataOut251) 
	 ,.R_out(R252) ,.data_out(dataOut252)  );
medianFilterCell  m253(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R252) ,.dataR_in(dataOut254) ,.dataL_in(dataOut252) 
	 ,.R_out(R253) ,.data_out(dataOut253)  );
medianFilterCell  m254(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R253) ,.dataR_in(dataOut255) ,.dataL_in(dataOut253) 
	 ,.R_out(R254) ,.data_out(dataOut254)  );
medianFilterCell  m255(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R254) ,.dataR_in(dataOut256) ,.dataL_in(dataOut254) 
	 ,.R_out(R255) ,.data_out(dataOut255)  );
medianFilterCell  m256(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R255) ,.dataR_in(dataOut257) ,.dataL_in(dataOut255) 
	 ,.R_out(R256) ,.data_out(dataOut256)  );
medianFilterCell  m257(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R256) ,.dataR_in(dataOut258) ,.dataL_in(dataOut256) 
	 ,.R_out(R257) ,.data_out(dataOut257)  );
medianFilterCell  m258(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R257) ,.dataR_in(dataOut259) ,.dataL_in(dataOut257) 
	 ,.R_out(R258) ,.data_out(dataOut258)  );
medianFilterCell  m259(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R258) ,.dataR_in(dataOut260) ,.dataL_in(dataOut258) 
	 ,.R_out(R259) ,.data_out(dataOut259)  );
medianFilterCell  m260(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R259) ,.dataR_in(dataOut261) ,.dataL_in(dataOut259) 
	 ,.R_out(R260) ,.data_out(dataOut260)  );
medianFilterCell  m261(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R260) ,.dataR_in(dataOut262) ,.dataL_in(dataOut260) 
	 ,.R_out(R261) ,.data_out(dataOut261)  );
medianFilterCell  m262(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R261) ,.dataR_in(dataOut263) ,.dataL_in(dataOut261) 
	 ,.R_out(R262) ,.data_out(dataOut262)  );
medianFilterCell  m263(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R262) ,.dataR_in(dataOut264) ,.dataL_in(dataOut262) 
	 ,.R_out(R263) ,.data_out(dataOut263)  );
medianFilterCell  m264(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R263) ,.dataR_in(dataOut265) ,.dataL_in(dataOut263) 
	 ,.R_out(R264) ,.data_out(dataOut264)  );
medianFilterCell  m265(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R264) ,.dataR_in(dataOut266) ,.dataL_in(dataOut264) 
	 ,.R_out(R265) ,.data_out(dataOut265)  );
medianFilterCell  m266(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R265) ,.dataR_in(dataOut267) ,.dataL_in(dataOut265) 
	 ,.R_out(R266) ,.data_out(dataOut266)  );
medianFilterCell  m267(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R266) ,.dataR_in(dataOut268) ,.dataL_in(dataOut266) 
	 ,.R_out(R267) ,.data_out(dataOut267)  );
medianFilterCell  m268(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R267) ,.dataR_in(dataOut269) ,.dataL_in(dataOut267) 
	 ,.R_out(R268) ,.data_out(dataOut268)  );
medianFilterCell  m269(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R268) ,.dataR_in(dataOut270) ,.dataL_in(dataOut268) 
	 ,.R_out(R269) ,.data_out(dataOut269)  );
medianFilterCell  m270(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R269) ,.dataR_in(dataOut271) ,.dataL_in(dataOut269) 
	 ,.R_out(R270) ,.data_out(dataOut270)  );
medianFilterCell  m271(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R270) ,.dataR_in(dataOut272) ,.dataL_in(dataOut270) 
	 ,.R_out(R271) ,.data_out(dataOut271)  );
medianFilterCell  m272(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R271) ,.dataR_in(dataOut273) ,.dataL_in(dataOut271) 
	 ,.R_out(R272) ,.data_out(dataOut272)  );
medianFilterCell  m273(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R272) ,.dataR_in(dataOut274) ,.dataL_in(dataOut272) 
	 ,.R_out(R273) ,.data_out(dataOut273)  );
medianFilterCell  m274(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R273) ,.dataR_in(dataOut275) ,.dataL_in(dataOut273) 
	 ,.R_out(R274) ,.data_out(dataOut274)  );
medianFilterCell  m275(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R274) ,.dataR_in(dataOut276) ,.dataL_in(dataOut274) 
	 ,.R_out(R275) ,.data_out(dataOut275)  );
medianFilterCell  m276(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R275) ,.dataR_in(dataOut277) ,.dataL_in(dataOut275) 
	 ,.R_out(R276) ,.data_out(dataOut276)  );
medianFilterCell  m277(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R276) ,.dataR_in(dataOut278) ,.dataL_in(dataOut276) 
	 ,.R_out(R277) ,.data_out(dataOut277)  );
medianFilterCell  m278(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R277) ,.dataR_in(dataOut279) ,.dataL_in(dataOut277) 
	 ,.R_out(R278) ,.data_out(dataOut278)  );
medianFilterCell  m279(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R278) ,.dataR_in(dataOut280) ,.dataL_in(dataOut278) 
	 ,.R_out(R279) ,.data_out(dataOut279)  );
medianFilterCell  m280(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R279) ,.dataR_in(dataOut281) ,.dataL_in(dataOut279) 
	 ,.R_out(R280) ,.data_out(dataOut280)  );
medianFilterCell  m281(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R280) ,.dataR_in(dataOut282) ,.dataL_in(dataOut280) 
	 ,.R_out(R281) ,.data_out(dataOut281)  );
medianFilterCell  m282(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R281) ,.dataR_in(dataOut283) ,.dataL_in(dataOut281) 
	 ,.R_out(R282) ,.data_out(dataOut282)  );
medianFilterCell  m283(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R282) ,.dataR_in(dataOut284) ,.dataL_in(dataOut282) 
	 ,.R_out(R283) ,.data_out(dataOut283)  );
medianFilterCell  m284(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R283) ,.dataR_in(dataOut285) ,.dataL_in(dataOut283) 
	 ,.R_out(R284) ,.data_out(dataOut284)  );
medianFilterCell  m285(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R284) ,.dataR_in(dataOut286) ,.dataL_in(dataOut284) 
	 ,.R_out(R285) ,.data_out(dataOut285)  );
medianFilterCell  m286(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R285) ,.dataR_in(dataOut287) ,.dataL_in(dataOut285) 
	 ,.R_out(R286) ,.data_out(dataOut286)  );
medianFilterCell  m287(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R286) ,.dataR_in(dataOut288) ,.dataL_in(dataOut286) 
	 ,.R_out(R287) ,.data_out(dataOut287)  );
medianFilterCell  m288(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R287) ,.dataR_in(dataOut289) ,.dataL_in(dataOut287) 
	 ,.R_out(R288) ,.data_out(dataOut288)  );
medianFilterCell  m289(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R288) ,.dataR_in(dataOut290) ,.dataL_in(dataOut288) 
	 ,.R_out(R289) ,.data_out(dataOut289)  );
medianFilterCell  m290(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R289) ,.dataR_in(dataOut291) ,.dataL_in(dataOut289) 
	 ,.R_out(R290) ,.data_out(dataOut290)  );
medianFilterCell  m291(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R290) ,.dataR_in(dataOut292) ,.dataL_in(dataOut290) 
	 ,.R_out(R291) ,.data_out(dataOut291)  );
medianFilterCell  m292(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R291) ,.dataR_in(dataOut293) ,.dataL_in(dataOut291) 
	 ,.R_out(R292) ,.data_out(dataOut292)  );
medianFilterCell  m293(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R292) ,.dataR_in(dataOut294) ,.dataL_in(dataOut292) 
	 ,.R_out(R293) ,.data_out(dataOut293)  );
medianFilterCell  m294(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R293) ,.dataR_in(dataOut295) ,.dataL_in(dataOut293) 
	 ,.R_out(R294) ,.data_out(dataOut294)  );
medianFilterCell  m295(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R294) ,.dataR_in(dataOut296) ,.dataL_in(dataOut294) 
	 ,.R_out(R295) ,.data_out(dataOut295)  );
medianFilterCell  m296(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R295) ,.dataR_in(dataOut297) ,.dataL_in(dataOut295) 
	 ,.R_out(R296) ,.data_out(dataOut296)  );
medianFilterCell  m297(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R296) ,.dataR_in(dataOut298) ,.dataL_in(dataOut296) 
	 ,.R_out(R297) ,.data_out(dataOut297)  );
medianFilterCell  m298(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R297) ,.dataR_in(dataOut299) ,.dataL_in(dataOut297) 
	 ,.R_out(R298) ,.data_out(dataOut298)  );
medianFilterCell  m299(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R298) ,.dataR_in(dataOut300) ,.dataL_in(dataOut298) 
	 ,.R_out(R299) ,.data_out(dataOut299)  );
medianFilterCell  m300(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R299) ,.dataR_in(dataOut301) ,.dataL_in(dataOut299) 
	 ,.R_out(R300) ,.data_out(dataOut300)  );
medianFilterCell  m301(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R300) ,.dataR_in(dataOut302) ,.dataL_in(dataOut300) 
	 ,.R_out(R301) ,.data_out(dataOut301)  );
medianFilterCell  m302(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R301) ,.dataR_in(dataOut303) ,.dataL_in(dataOut301) 
	 ,.R_out(R302) ,.data_out(dataOut302)  );
medianFilterCell  m303(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R302) ,.dataR_in(dataOut304) ,.dataL_in(dataOut302) 
	 ,.R_out(R303) ,.data_out(dataOut303)  );
medianFilterCell  m304(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R303) ,.dataR_in(dataOut305) ,.dataL_in(dataOut303) 
	 ,.R_out(R304) ,.data_out(dataOut304)  );
medianFilterCell  m305(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R304) ,.dataR_in(dataOut306) ,.dataL_in(dataOut304) 
	 ,.R_out(R305) ,.data_out(dataOut305)  );
medianFilterCell  m306(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R305) ,.dataR_in(dataOut307) ,.dataL_in(dataOut305) 
	 ,.R_out(R306) ,.data_out(dataOut306)  );
medianFilterCell  m307(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R306) ,.dataR_in(dataOut308) ,.dataL_in(dataOut306) 
	 ,.R_out(R307) ,.data_out(dataOut307)  );
medianFilterCell  m308(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R307) ,.dataR_in(dataOut309) ,.dataL_in(dataOut307) 
	 ,.R_out(R308) ,.data_out(dataOut308)  );
medianFilterCell  m309(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R308) ,.dataR_in(dataOut310) ,.dataL_in(dataOut308) 
	 ,.R_out(R309) ,.data_out(dataOut309)  );
medianFilterCell  m310(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R309) ,.dataR_in(dataOut311) ,.dataL_in(dataOut309) 
	 ,.R_out(R310) ,.data_out(dataOut310)  );
medianFilterCell  m311(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R310) ,.dataR_in(dataOut312) ,.dataL_in(dataOut310) 
	 ,.R_out(R311) ,.data_out(dataOut311)  );
medianFilterCell  m312(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R311) ,.dataR_in(dataOut313) ,.dataL_in(dataOut311) 
	 ,.R_out(R312) ,.data_out(dataOut312)  );
medianFilterCell  m313(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R312) ,.dataR_in(dataOut314) ,.dataL_in(dataOut312) 
	 ,.R_out(R313) ,.data_out(dataOut313)  );
medianFilterCell  m314(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R313) ,.dataR_in(dataOut315) ,.dataL_in(dataOut313) 
	 ,.R_out(R314) ,.data_out(dataOut314)  );
medianFilterCell  m315(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R314) ,.dataR_in(dataOut316) ,.dataL_in(dataOut314) 
	 ,.R_out(R315) ,.data_out(dataOut315)  );
medianFilterCell  m316(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R315) ,.dataR_in(dataOut317) ,.dataL_in(dataOut315) 
	 ,.R_out(R316) ,.data_out(dataOut316)  );
medianFilterCell  m317(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R316) ,.dataR_in(dataOut318) ,.dataL_in(dataOut316) 
	 ,.R_out(R317) ,.data_out(dataOut317)  );
medianFilterCell  m318(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R317) ,.dataR_in(dataOut319) ,.dataL_in(dataOut317) 
	 ,.R_out(R318) ,.data_out(dataOut318)  );
medianFilterCell  m319(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R318) ,.dataR_in(dataOut320) ,.dataL_in(dataOut318) 
	 ,.R_out(R319) ,.data_out(dataOut319)  );
medianFilterCell  m320(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R319) ,.dataR_in(dataOut321) ,.dataL_in(dataOut319) 
	 ,.R_out(R320) ,.data_out(dataOut320)  );
medianFilterCell  m321(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R320) ,.dataR_in(dataOut322) ,.dataL_in(dataOut320) 
	 ,.R_out(R321) ,.data_out(dataOut321)  );
medianFilterCell  m322(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R321) ,.dataR_in(dataOut323) ,.dataL_in(dataOut321) 
	 ,.R_out(R322) ,.data_out(dataOut322)  );
medianFilterCell  m323(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R322) ,.dataR_in(dataOut324) ,.dataL_in(dataOut322) 
	 ,.R_out(R323) ,.data_out(dataOut323)  );
medianFilterCell  m324(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R323) ,.dataR_in(dataOut325) ,.dataL_in(dataOut323) 
	 ,.R_out(R324) ,.data_out(dataOut324)  );
medianFilterCell  m325(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R324) ,.dataR_in(dataOut326) ,.dataL_in(dataOut324) 
	 ,.R_out(R325) ,.data_out(dataOut325)  );
medianFilterCell  m326(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R325) ,.dataR_in(dataOut327) ,.dataL_in(dataOut325) 
	 ,.R_out(R326) ,.data_out(dataOut326)  );
medianFilterCell  m327(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R326) ,.dataR_in(dataOut328) ,.dataL_in(dataOut326) 
	 ,.R_out(R327) ,.data_out(dataOut327)  );
medianFilterCell  m328(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R327) ,.dataR_in(dataOut329) ,.dataL_in(dataOut327) 
	 ,.R_out(R328) ,.data_out(dataOut328)  );
medianFilterCell  m329(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R328) ,.dataR_in(dataOut330) ,.dataL_in(dataOut328) 
	 ,.R_out(R329) ,.data_out(dataOut329)  );
medianFilterCell  m330(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R329) ,.dataR_in(dataOut331) ,.dataL_in(dataOut329) 
	 ,.R_out(R330) ,.data_out(dataOut330)  );
medianFilterCell  m331(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R330) ,.dataR_in(dataOut332) ,.dataL_in(dataOut330) 
	 ,.R_out(R331) ,.data_out(dataOut331)  );
medianFilterCell  m332(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R331) ,.dataR_in(dataOut333) ,.dataL_in(dataOut331) 
	 ,.R_out(R332) ,.data_out(dataOut332)  );
medianFilterCell  m333(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R332) ,.dataR_in(dataOut334) ,.dataL_in(dataOut332) 
	 ,.R_out(R333) ,.data_out(dataOut333)  );
medianFilterCell  m334(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R333) ,.dataR_in(dataOut335) ,.dataL_in(dataOut333) 
	 ,.R_out(R334) ,.data_out(dataOut334)  );
medianFilterCell  m335(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R334) ,.dataR_in(dataOut336) ,.dataL_in(dataOut334) 
	 ,.R_out(R335) ,.data_out(dataOut335)  );
medianFilterCell  m336(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R335) ,.dataR_in(dataOut337) ,.dataL_in(dataOut335) 
	 ,.R_out(R336) ,.data_out(dataOut336)  );
medianFilterCell  m337(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R336) ,.dataR_in(dataOut338) ,.dataL_in(dataOut336) 
	 ,.R_out(R337) ,.data_out(dataOut337)  );
medianFilterCell  m338(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R337) ,.dataR_in(dataOut339) ,.dataL_in(dataOut337) 
	 ,.R_out(R338) ,.data_out(dataOut338)  );
medianFilterCell  m339(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R338) ,.dataR_in(dataOut340) ,.dataL_in(dataOut338) 
	 ,.R_out(R339) ,.data_out(dataOut339)  );
medianFilterCell  m340(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R339) ,.dataR_in(dataOut341) ,.dataL_in(dataOut339) 
	 ,.R_out(R340) ,.data_out(dataOut340)  );
medianFilterCell  m341(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R340) ,.dataR_in(dataOut342) ,.dataL_in(dataOut340) 
	 ,.R_out(R341) ,.data_out(dataOut341)  );
medianFilterCell  m342(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R341) ,.dataR_in(dataOut343) ,.dataL_in(dataOut341) 
	 ,.R_out(R342) ,.data_out(dataOut342)  );
medianFilterCell  m343(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R342) ,.dataR_in(dataOut344) ,.dataL_in(dataOut342) 
	 ,.R_out(R343) ,.data_out(dataOut343)  );
medianFilterCell  m344(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R343) ,.dataR_in(dataOut345) ,.dataL_in(dataOut343) 
	 ,.R_out(R344) ,.data_out(dataOut344)  );
medianFilterCell  m345(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R344) ,.dataR_in(dataOut346) ,.dataL_in(dataOut344) 
	 ,.R_out(R345) ,.data_out(dataOut345)  );
medianFilterCell  m346(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R345) ,.dataR_in(dataOut347) ,.dataL_in(dataOut345) 
	 ,.R_out(R346) ,.data_out(dataOut346)  );
medianFilterCell  m347(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R346) ,.dataR_in(dataOut348) ,.dataL_in(dataOut346) 
	 ,.R_out(R347) ,.data_out(dataOut347)  );
medianFilterCell  m348(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R347) ,.dataR_in(dataOut349) ,.dataL_in(dataOut347) 
	 ,.R_out(R348) ,.data_out(dataOut348)  );
medianFilterCell  m349(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R348) ,.dataR_in(dataOut350) ,.dataL_in(dataOut348) 
	 ,.R_out(R349) ,.data_out(dataOut349)  );
medianFilterCell  m350(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R349) ,.dataR_in(dataOut351) ,.dataL_in(dataOut349) 
	 ,.R_out(R350) ,.data_out(dataOut350)  );
medianFilterCell  m351(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R350) ,.dataR_in(dataOut352) ,.dataL_in(dataOut350) 
	 ,.R_out(R351) ,.data_out(dataOut351)  );
medianFilterCell  m352(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R351) ,.dataR_in(dataOut353) ,.dataL_in(dataOut351) 
	 ,.R_out(R352) ,.data_out(dataOut352)  );
medianFilterCell  m353(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R352) ,.dataR_in(dataOut354) ,.dataL_in(dataOut352) 
	 ,.R_out(R353) ,.data_out(dataOut353)  );
medianFilterCell  m354(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R353) ,.dataR_in(dataOut355) ,.dataL_in(dataOut353) 
	 ,.R_out(R354) ,.data_out(dataOut354)  );
medianFilterCell  m355(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R354) ,.dataR_in(dataOut356) ,.dataL_in(dataOut354) 
	 ,.R_out(R355) ,.data_out(dataOut355)  );
medianFilterCell  m356(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R355) ,.dataR_in(dataOut357) ,.dataL_in(dataOut355) 
	 ,.R_out(R356) ,.data_out(dataOut356)  );
medianFilterCell  m357(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R356) ,.dataR_in(dataOut358) ,.dataL_in(dataOut356) 
	 ,.R_out(R357) ,.data_out(dataOut357)  );
medianFilterCell  m358(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R357) ,.dataR_in(dataOut359) ,.dataL_in(dataOut357) 
	 ,.R_out(R358) ,.data_out(dataOut358)  );
medianFilterCell  m359(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R358) ,.dataR_in(dataOut360) ,.dataL_in(dataOut358) 
	 ,.R_out(R359) ,.data_out(dataOut359)  );
medianFilterCell  m360(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R359) ,.dataR_in(dataOut361) ,.dataL_in(dataOut359) 
	 ,.R_out(R360) ,.data_out(dataOut360)  );
medianFilterCell  m361(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R360) ,.dataR_in(dataOut362) ,.dataL_in(dataOut360) 
	 ,.R_out(R361) ,.data_out(dataOut361)  );
medianFilterCell  m362(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R361) ,.dataR_in(dataOut363) ,.dataL_in(dataOut361) 
	 ,.R_out(R362) ,.data_out(dataOut362)  );
medianFilterCell  m363(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R362) ,.dataR_in(dataOut364) ,.dataL_in(dataOut362) 
	 ,.R_out(R363) ,.data_out(dataOut363)  );
medianFilterCell  m364(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R363) ,.dataR_in(dataOut365) ,.dataL_in(dataOut363) 
	 ,.R_out(R364) ,.data_out(dataOut364)  );
medianFilterCell  m365(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R364) ,.dataR_in(dataOut366) ,.dataL_in(dataOut364) 
	 ,.R_out(R365) ,.data_out(dataOut365)  );
medianFilterCell  m366(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R365) ,.dataR_in(dataOut367) ,.dataL_in(dataOut365) 
	 ,.R_out(R366) ,.data_out(dataOut366)  );
medianFilterCell  m367(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R366) ,.dataR_in(dataOut368) ,.dataL_in(dataOut366) 
	 ,.R_out(R367) ,.data_out(dataOut367)  );
medianFilterCell  m368(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R367) ,.dataR_in(dataOut369) ,.dataL_in(dataOut367) 
	 ,.R_out(R368) ,.data_out(dataOut368)  );
medianFilterCell  m369(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R368) ,.dataR_in(dataOut370) ,.dataL_in(dataOut368) 
	 ,.R_out(R369) ,.data_out(dataOut369)  );
medianFilterCell  m370(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R369) ,.dataR_in(dataOut371) ,.dataL_in(dataOut369) 
	 ,.R_out(R370) ,.data_out(dataOut370)  );
medianFilterCell  m371(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R370) ,.dataR_in(dataOut372) ,.dataL_in(dataOut370) 
	 ,.R_out(R371) ,.data_out(dataOut371)  );
medianFilterCell  m372(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R371) ,.dataR_in(dataOut373) ,.dataL_in(dataOut371) 
	 ,.R_out(R372) ,.data_out(dataOut372)  );
medianFilterCell  m373(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R372) ,.dataR_in(dataOut374) ,.dataL_in(dataOut372) 
	 ,.R_out(R373) ,.data_out(dataOut373)  );
medianFilterCell  m374(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R373) ,.dataR_in(dataOut375) ,.dataL_in(dataOut373) 
	 ,.R_out(R374) ,.data_out(dataOut374)  );
medianFilterCell  m375(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R374) ,.dataR_in(dataOut376) ,.dataL_in(dataOut374) 
	 ,.R_out(R375) ,.data_out(dataOut375)  );
medianFilterCell  m376(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R375) ,.dataR_in(dataOut377) ,.dataL_in(dataOut375) 
	 ,.R_out(R376) ,.data_out(dataOut376)  );
medianFilterCell  m377(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R376) ,.dataR_in(dataOut378) ,.dataL_in(dataOut376) 
	 ,.R_out(R377) ,.data_out(dataOut377)  );
medianFilterCell  m378(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R377) ,.dataR_in(dataOut379) ,.dataL_in(dataOut377) 
	 ,.R_out(R378) ,.data_out(dataOut378)  );
medianFilterCell  m379(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R378) ,.dataR_in(dataOut380) ,.dataL_in(dataOut378) 
	 ,.R_out(R379) ,.data_out(dataOut379)  );
medianFilterCell  m380(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R379) ,.dataR_in(dataOut381) ,.dataL_in(dataOut379) 
	 ,.R_out(R380) ,.data_out(dataOut380)  );
medianFilterCell  m381(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R380) ,.dataR_in(dataOut382) ,.dataL_in(dataOut380) 
	 ,.R_out(R381) ,.data_out(dataOut381)  );
medianFilterCell  m382(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R381) ,.dataR_in(dataOut383) ,.dataL_in(dataOut381) 
	 ,.R_out(R382) ,.data_out(dataOut382)  );
medianFilterCell  m383(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R382) ,.dataR_in(dataOut384) ,.dataL_in(dataOut382) 
	 ,.R_out(R383) ,.data_out(dataOut383)  );
medianFilterCell  m384(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R383) ,.dataR_in(dataOut385) ,.dataL_in(dataOut383) 
	 ,.R_out(R384) ,.data_out(dataOut384)  );
medianFilterCell  m385(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R384) ,.dataR_in(dataOut386) ,.dataL_in(dataOut384) 
	 ,.R_out(R385) ,.data_out(dataOut385)  );
medianFilterCell  m386(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R385) ,.dataR_in(dataOut387) ,.dataL_in(dataOut385) 
	 ,.R_out(R386) ,.data_out(dataOut386)  );
medianFilterCell  m387(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R386) ,.dataR_in(dataOut388) ,.dataL_in(dataOut386) 
	 ,.R_out(R387) ,.data_out(dataOut387)  );
medianFilterCell  m388(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R387) ,.dataR_in(dataOut389) ,.dataL_in(dataOut387) 
	 ,.R_out(R388) ,.data_out(dataOut388)  );
medianFilterCell  m389(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R388) ,.dataR_in(dataOut390) ,.dataL_in(dataOut388) 
	 ,.R_out(R389) ,.data_out(dataOut389)  );
medianFilterCell  m390(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R389) ,.dataR_in(dataOut391) ,.dataL_in(dataOut389) 
	 ,.R_out(R390) ,.data_out(dataOut390)  );
medianFilterCell  m391(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R390) ,.dataR_in(dataOut392) ,.dataL_in(dataOut390) 
	 ,.R_out(R391) ,.data_out(dataOut391)  );
medianFilterCell  m392(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R391) ,.dataR_in(dataOut393) ,.dataL_in(dataOut391) 
	 ,.R_out(R392) ,.data_out(dataOut392)  );
medianFilterCell  m393(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R392) ,.dataR_in(dataOut394) ,.dataL_in(dataOut392) 
	 ,.R_out(R393) ,.data_out(dataOut393)  );
medianFilterCell  m394(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R393) ,.dataR_in(dataOut395) ,.dataL_in(dataOut393) 
	 ,.R_out(R394) ,.data_out(dataOut394)  );
medianFilterCell  m395(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R394) ,.dataR_in(dataOut396) ,.dataL_in(dataOut394) 
	 ,.R_out(R395) ,.data_out(dataOut395)  );
medianFilterCell  m396(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R395) ,.dataR_in(dataOut397) ,.dataL_in(dataOut395) 
	 ,.R_out(R396) ,.data_out(dataOut396)  );
medianFilterCell  m397(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R396) ,.dataR_in(dataOut398) ,.dataL_in(dataOut396) 
	 ,.R_out(R397) ,.data_out(dataOut397)  );
medianFilterCell  m398(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R397) ,.dataR_in(dataOut399) ,.dataL_in(dataOut397) 
	 ,.R_out(R398) ,.data_out(dataOut398)  );
medianFilterCell  m399(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R398) ,.dataR_in(dataOut400) ,.dataL_in(dataOut398) 
	 ,.R_out(R399) ,.data_out(dataOut399)  );
medianFilterCell  m400(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R399) ,.dataR_in(dataOut401) ,.dataL_in(dataOut399) 
	 ,.R_out(R400) ,.data_out(dataOut400)  );
medianFilterCell  m401(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R400) ,.dataR_in(dataOut402) ,.dataL_in(dataOut400) 
	 ,.R_out(R401) ,.data_out(dataOut401)  );
medianFilterCell  m402(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R401) ,.dataR_in(dataOut403) ,.dataL_in(dataOut401) 
	 ,.R_out(R402) ,.data_out(dataOut402)  );
medianFilterCell  m403(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R402) ,.dataR_in(dataOut404) ,.dataL_in(dataOut402) 
	 ,.R_out(R403) ,.data_out(dataOut403)  );
medianFilterCell  m404(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R403) ,.dataR_in(dataOut405) ,.dataL_in(dataOut403) 
	 ,.R_out(R404) ,.data_out(dataOut404)  );
medianFilterCell  m405(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R404) ,.dataR_in(dataOut406) ,.dataL_in(dataOut404) 
	 ,.R_out(R405) ,.data_out(dataOut405)  );
medianFilterCell  m406(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R405) ,.dataR_in(dataOut407) ,.dataL_in(dataOut405) 
	 ,.R_out(R406) ,.data_out(dataOut406)  );
medianFilterCell  m407(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R406) ,.dataR_in(dataOut408) ,.dataL_in(dataOut406) 
	 ,.R_out(R407) ,.data_out(dataOut407)  );
medianFilterCell  m408(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R407) ,.dataR_in(dataOut409) ,.dataL_in(dataOut407) 
	 ,.R_out(R408) ,.data_out(dataOut408)  );
medianFilterCell  m409(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R408) ,.dataR_in(dataOut410) ,.dataL_in(dataOut408) 
	 ,.R_out(R409) ,.data_out(dataOut409)  );
medianFilterCell  m410(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R409) ,.dataR_in(dataOut411) ,.dataL_in(dataOut409) 
	 ,.R_out(R410) ,.data_out(dataOut410)  );
medianFilterCell  m411(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R410) ,.dataR_in(dataOut412) ,.dataL_in(dataOut410) 
	 ,.R_out(R411) ,.data_out(dataOut411)  );
medianFilterCell  m412(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R411) ,.dataR_in(dataOut413) ,.dataL_in(dataOut411) 
	 ,.R_out(R412) ,.data_out(dataOut412)  );
medianFilterCell  m413(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R412) ,.dataR_in(dataOut414) ,.dataL_in(dataOut412) 
	 ,.R_out(R413) ,.data_out(dataOut413)  );
medianFilterCell  m414(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R413) ,.dataR_in(dataOut415) ,.dataL_in(dataOut413) 
	 ,.R_out(R414) ,.data_out(dataOut414)  );
medianFilterCell  m415(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R414) ,.dataR_in(dataOut416) ,.dataL_in(dataOut414) 
	 ,.R_out(R415) ,.data_out(dataOut415)  );
medianFilterCell  m416(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R415) ,.dataR_in(dataOut417) ,.dataL_in(dataOut415) 
	 ,.R_out(R416) ,.data_out(dataOut416)  );
medianFilterCell  m417(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R416) ,.dataR_in(dataOut418) ,.dataL_in(dataOut416) 
	 ,.R_out(R417) ,.data_out(dataOut417)  );
medianFilterCell  m418(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R417) ,.dataR_in(dataOut419) ,.dataL_in(dataOut417) 
	 ,.R_out(R418) ,.data_out(dataOut418)  );
medianFilterCell  m419(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R418) ,.dataR_in(dataOut420) ,.dataL_in(dataOut418) 
	 ,.R_out(R419) ,.data_out(dataOut419)  );
medianFilterCell  m420(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R419) ,.dataR_in(dataOut421) ,.dataL_in(dataOut419) 
	 ,.R_out(R420) ,.data_out(dataOut420)  );
medianFilterCell  m421(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R420) ,.dataR_in(dataOut422) ,.dataL_in(dataOut420) 
	 ,.R_out(R421) ,.data_out(dataOut421)  );
medianFilterCell  m422(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R421) ,.dataR_in(dataOut423) ,.dataL_in(dataOut421) 
	 ,.R_out(R422) ,.data_out(dataOut422)  );
medianFilterCell  m423(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R422) ,.dataR_in(dataOut424) ,.dataL_in(dataOut422) 
	 ,.R_out(R423) ,.data_out(dataOut423)  );
medianFilterCell  m424(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R423) ,.dataR_in(dataOut425) ,.dataL_in(dataOut423) 
	 ,.R_out(R424) ,.data_out(dataOut424)  );
medianFilterCell  m425(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R424) ,.dataR_in(dataOut426) ,.dataL_in(dataOut424) 
	 ,.R_out(R425) ,.data_out(dataOut425)  );
medianFilterCell  m426(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R425) ,.dataR_in(dataOut427) ,.dataL_in(dataOut425) 
	 ,.R_out(R426) ,.data_out(dataOut426)  );
medianFilterCell  m427(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R426) ,.dataR_in(dataOut428) ,.dataL_in(dataOut426) 
	 ,.R_out(R427) ,.data_out(dataOut427)  );
medianFilterCell  m428(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R427) ,.dataR_in(dataOut429) ,.dataL_in(dataOut427) 
	 ,.R_out(R428) ,.data_out(dataOut428)  );
medianFilterCell  m429(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R428) ,.dataR_in(dataOut430) ,.dataL_in(dataOut428) 
	 ,.R_out(R429) ,.data_out(dataOut429)  );
medianFilterCell  m430(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R429) ,.dataR_in(dataOut431) ,.dataL_in(dataOut429) 
	 ,.R_out(R430) ,.data_out(dataOut430)  );
medianFilterCell  m431(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R430) ,.dataR_in(dataOut432) ,.dataL_in(dataOut430) 
	 ,.R_out(R431) ,.data_out(dataOut431)  );
medianFilterCell  m432(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R431) ,.dataR_in(dataOut433) ,.dataL_in(dataOut431) 
	 ,.R_out(R432) ,.data_out(dataOut432)  );
medianFilterCell  m433(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R432) ,.dataR_in(dataOut434) ,.dataL_in(dataOut432) 
	 ,.R_out(R433) ,.data_out(dataOut433)  );
medianFilterCell  m434(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R433) ,.dataR_in(dataOut435) ,.dataL_in(dataOut433) 
	 ,.R_out(R434) ,.data_out(dataOut434)  );
medianFilterCell  m435(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R434) ,.dataR_in(dataOut436) ,.dataL_in(dataOut434) 
	 ,.R_out(R435) ,.data_out(dataOut435)  );
medianFilterCell  m436(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R435) ,.dataR_in(dataOut437) ,.dataL_in(dataOut435) 
	 ,.R_out(R436) ,.data_out(dataOut436)  );
medianFilterCell  m437(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R436) ,.dataR_in(dataOut438) ,.dataL_in(dataOut436) 
	 ,.R_out(R437) ,.data_out(dataOut437)  );
medianFilterCell  m438(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R437) ,.dataR_in(dataOut439) ,.dataL_in(dataOut437) 
	 ,.R_out(R438) ,.data_out(dataOut438)  );
medianFilterCell  m439(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R438) ,.dataR_in(dataOut440) ,.dataL_in(dataOut438) 
	 ,.R_out(R439) ,.data_out(dataOut439)  );
medianFilterCell  m440(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R439) ,.dataR_in(dataOut441) ,.dataL_in(dataOut439) 
	 ,.R_out(R440) ,.data_out(dataOut440)  );
medianFilterCell  m441(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R440) ,.dataR_in(dataOut442) ,.dataL_in(dataOut440) 
	 ,.R_out(R441) ,.data_out(dataOut441)  );
medianFilterCell  m442(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R441) ,.dataR_in(dataOut443) ,.dataL_in(dataOut441) 
	 ,.R_out(R442) ,.data_out(dataOut442)  );
medianFilterCell  m443(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R442) ,.dataR_in(dataOut444) ,.dataL_in(dataOut442) 
	 ,.R_out(R443) ,.data_out(dataOut443)  );
medianFilterCell  m444(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R443) ,.dataR_in(dataOut445) ,.dataL_in(dataOut443) 
	 ,.R_out(R444) ,.data_out(dataOut444)  );
medianFilterCell  m445(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R444) ,.dataR_in(dataOut446) ,.dataL_in(dataOut444) 
	 ,.R_out(R445) ,.data_out(dataOut445)  );
medianFilterCell  m446(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R445) ,.dataR_in(dataOut447) ,.dataL_in(dataOut445) 
	 ,.R_out(R446) ,.data_out(dataOut446)  );
medianFilterCell  m447(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R446) ,.dataR_in(dataOut448) ,.dataL_in(dataOut446) 
	 ,.R_out(R447) ,.data_out(dataOut447)  );
medianFilterCell  m448(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R447) ,.dataR_in(dataOut449) ,.dataL_in(dataOut447) 
	 ,.R_out(R448) ,.data_out(dataOut448)  );
medianFilterCell  m449(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R448) ,.dataR_in(dataOut450) ,.dataL_in(dataOut448) 
	 ,.R_out(R449) ,.data_out(dataOut449)  );
medianFilterCell  m450(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R449) ,.dataR_in(dataOut451) ,.dataL_in(dataOut449) 
	 ,.R_out(R450) ,.data_out(dataOut450)  );
medianFilterCell  m451(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R450) ,.dataR_in(dataOut452) ,.dataL_in(dataOut450) 
	 ,.R_out(R451) ,.data_out(dataOut451)  );
medianFilterCell  m452(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R451) ,.dataR_in(dataOut453) ,.dataL_in(dataOut451) 
	 ,.R_out(R452) ,.data_out(dataOut452)  );
medianFilterCell  m453(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R452) ,.dataR_in(dataOut454) ,.dataL_in(dataOut452) 
	 ,.R_out(R453) ,.data_out(dataOut453)  );
medianFilterCell  m454(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R453) ,.dataR_in(dataOut455) ,.dataL_in(dataOut453) 
	 ,.R_out(R454) ,.data_out(dataOut454)  );
medianFilterCell  m455(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R454) ,.dataR_in(dataOut456) ,.dataL_in(dataOut454) 
	 ,.R_out(R455) ,.data_out(dataOut455)  );
medianFilterCell  m456(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R455) ,.dataR_in(dataOut457) ,.dataL_in(dataOut455) 
	 ,.R_out(R456) ,.data_out(dataOut456)  );
medianFilterCell  m457(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R456) ,.dataR_in(dataOut458) ,.dataL_in(dataOut456) 
	 ,.R_out(R457) ,.data_out(dataOut457)  );
medianFilterCell  m458(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R457) ,.dataR_in(dataOut459) ,.dataL_in(dataOut457) 
	 ,.R_out(R458) ,.data_out(dataOut458)  );
medianFilterCell  m459(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R458) ,.dataR_in(dataOut460) ,.dataL_in(dataOut458) 
	 ,.R_out(R459) ,.data_out(dataOut459)  );
medianFilterCell  m460(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R459) ,.dataR_in(dataOut461) ,.dataL_in(dataOut459) 
	 ,.R_out(R460) ,.data_out(dataOut460)  );
medianFilterCell  m461(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R460) ,.dataR_in(dataOut462) ,.dataL_in(dataOut460) 
	 ,.R_out(R461) ,.data_out(dataOut461)  );
medianFilterCell  m462(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R461) ,.dataR_in(dataOut463) ,.dataL_in(dataOut461) 
	 ,.R_out(R462) ,.data_out(dataOut462)  );
medianFilterCell  m463(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R462) ,.dataR_in(dataOut464) ,.dataL_in(dataOut462) 
	 ,.R_out(R463) ,.data_out(dataOut463)  );
medianFilterCell  m464(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R463) ,.dataR_in(dataOut465) ,.dataL_in(dataOut463) 
	 ,.R_out(R464) ,.data_out(dataOut464)  );
medianFilterCell  m465(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R464) ,.dataR_in(dataOut466) ,.dataL_in(dataOut464) 
	 ,.R_out(R465) ,.data_out(dataOut465)  );
medianFilterCell  m466(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R465) ,.dataR_in(dataOut467) ,.dataL_in(dataOut465) 
	 ,.R_out(R466) ,.data_out(dataOut466)  );
medianFilterCell  m467(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R466) ,.dataR_in(dataOut468) ,.dataL_in(dataOut466) 
	 ,.R_out(R467) ,.data_out(dataOut467)  );
medianFilterCell  m468(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R467) ,.dataR_in(dataOut469) ,.dataL_in(dataOut467) 
	 ,.R_out(R468) ,.data_out(dataOut468)  );
medianFilterCell  m469(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R468) ,.dataR_in(dataOut470) ,.dataL_in(dataOut468) 
	 ,.R_out(R469) ,.data_out(dataOut469)  );
medianFilterCell  m470(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R469) ,.dataR_in(dataOut471) ,.dataL_in(dataOut469) 
	 ,.R_out(R470) ,.data_out(dataOut470)  );
medianFilterCell  m471(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R470) ,.dataR_in(dataOut472) ,.dataL_in(dataOut470) 
	 ,.R_out(R471) ,.data_out(dataOut471)  );
medianFilterCell  m472(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R471) ,.dataR_in(dataOut473) ,.dataL_in(dataOut471) 
	 ,.R_out(R472) ,.data_out(dataOut472)  );
medianFilterCell  m473(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R472) ,.dataR_in(dataOut474) ,.dataL_in(dataOut472) 
	 ,.R_out(R473) ,.data_out(dataOut473)  );
medianFilterCell  m474(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R473) ,.dataR_in(dataOut475) ,.dataL_in(dataOut473) 
	 ,.R_out(R474) ,.data_out(dataOut474)  );
medianFilterCell  m475(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R474) ,.dataR_in(dataOut476) ,.dataL_in(dataOut474) 
	 ,.R_out(R475) ,.data_out(dataOut475)  );
medianFilterCell  m476(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R475) ,.dataR_in(dataOut477) ,.dataL_in(dataOut475) 
	 ,.R_out(R476) ,.data_out(dataOut476)  );
medianFilterCell  m477(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R476) ,.dataR_in(dataOut478) ,.dataL_in(dataOut476) 
	 ,.R_out(R477) ,.data_out(dataOut477)  );
medianFilterCell  m478(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R477) ,.dataR_in(dataOut479) ,.dataL_in(dataOut477) 
	 ,.R_out(R478) ,.data_out(dataOut478)  );
medianFilterCell  m479(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R478) ,.dataR_in(dataOut480) ,.dataL_in(dataOut478) 
	 ,.R_out(R479) ,.data_out(dataOut479)  );
medianFilterCell  m480(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R479) ,.dataR_in(dataOut481) ,.dataL_in(dataOut479) 
	 ,.R_out(R480) ,.data_out(dataOut480)  );
medianFilterCell  m481(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R480) ,.dataR_in(dataOut482) ,.dataL_in(dataOut480) 
	 ,.R_out(R481) ,.data_out(dataOut481)  );
medianFilterCell  m482(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R481) ,.dataR_in(dataOut483) ,.dataL_in(dataOut481) 
	 ,.R_out(R482) ,.data_out(dataOut482)  );
medianFilterCell  m483(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R482) ,.dataR_in(dataOut484) ,.dataL_in(dataOut482) 
	 ,.R_out(R483) ,.data_out(dataOut483)  );
medianFilterCell  m484(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R483) ,.dataR_in(dataOut485) ,.dataL_in(dataOut483) 
	 ,.R_out(R484) ,.data_out(dataOut484)  );
medianFilterCell  m485(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R484) ,.dataR_in(dataOut486) ,.dataL_in(dataOut484) 
	 ,.R_out(R485) ,.data_out(dataOut485)  );
medianFilterCell  m486(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R485) ,.dataR_in(dataOut487) ,.dataL_in(dataOut485) 
	 ,.R_out(R486) ,.data_out(dataOut486)  );
medianFilterCell  m487(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R486) ,.dataR_in(dataOut488) ,.dataL_in(dataOut486) 
	 ,.R_out(R487) ,.data_out(dataOut487)  );
medianFilterCell  m488(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R487) ,.dataR_in(dataOut489) ,.dataL_in(dataOut487) 
	 ,.R_out(R488) ,.data_out(dataOut488)  );
medianFilterCell  m489(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R488) ,.dataR_in(dataOut490) ,.dataL_in(dataOut488) 
	 ,.R_out(R489) ,.data_out(dataOut489)  );
medianFilterCell  m490(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R489) ,.dataR_in(dataOut491) ,.dataL_in(dataOut489) 
	 ,.R_out(R490) ,.data_out(dataOut490)  );
medianFilterCell  m491(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R490) ,.dataR_in(dataOut492) ,.dataL_in(dataOut490) 
	 ,.R_out(R491) ,.data_out(dataOut491)  );
medianFilterCell  m492(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R491) ,.dataR_in(dataOut493) ,.dataL_in(dataOut491) 
	 ,.R_out(R492) ,.data_out(dataOut492)  );
medianFilterCell  m493(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R492) ,.dataR_in(dataOut494) ,.dataL_in(dataOut492) 
	 ,.R_out(R493) ,.data_out(dataOut493)  );
medianFilterCell  m494(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R493) ,.dataR_in(dataOut495) ,.dataL_in(dataOut493) 
	 ,.R_out(R494) ,.data_out(dataOut494)  );
medianFilterCell  m495(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R494) ,.dataR_in(dataOut496) ,.dataL_in(dataOut494) 
	 ,.R_out(R495) ,.data_out(dataOut495)  );
medianFilterCell  m496(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R495) ,.dataR_in(dataOut497) ,.dataL_in(dataOut495) 
	 ,.R_out(R496) ,.data_out(dataOut496)  );
medianFilterCell  m497(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R496) ,.dataR_in(dataOut498) ,.dataL_in(dataOut496) 
	 ,.R_out(R497) ,.data_out(dataOut497)  );
medianFilterCell  m498(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R497) ,.dataR_in(dataOut499) ,.dataL_in(dataOut497) 
	 ,.R_out(R498) ,.data_out(dataOut498)  );
medianFilterCell  m499(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R498) ,.dataR_in(dataOut500) ,.dataL_in(dataOut498) 
	 ,.R_out(R499) ,.data_out(dataOut499)  );
medianFilterCell  m500(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R499) ,.dataR_in(dataOut501) ,.dataL_in(dataOut499) 
	 ,.R_out(R500) ,.data_out(dataOut500)  );
medianFilterCell  m501(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R500) ,.dataR_in(dataOut502) ,.dataL_in(dataOut500) 
	 ,.R_out(R501) ,.data_out(dataOut501)  );
medianFilterCell  m502(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R501) ,.dataR_in(dataOut503) ,.dataL_in(dataOut501) 
	 ,.R_out(R502) ,.data_out(dataOut502)  );
medianFilterCell  m503(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R502) ,.dataR_in(dataOut504) ,.dataL_in(dataOut502) 
	 ,.R_out(R503) ,.data_out(dataOut503)  );
medianFilterCell  m504(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R503) ,.dataR_in(dataOut505) ,.dataL_in(dataOut503) 
	 ,.R_out(R504) ,.data_out(dataOut504)  );
medianFilterCell  m505(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R504) ,.dataR_in(dataOut506) ,.dataL_in(dataOut504) 
	 ,.R_out(R505) ,.data_out(dataOut505)  );
medianFilterCell  m506(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R505) ,.dataR_in(dataOut507) ,.dataL_in(dataOut505) 
	 ,.R_out(R506) ,.data_out(dataOut506)  );
medianFilterCell  m507(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R506) ,.dataR_in(dataOut508) ,.dataL_in(dataOut506) 
	 ,.R_out(R507) ,.data_out(dataOut507)  );
medianFilterCell  m508(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R507) ,.dataR_in(dataOut509) ,.dataL_in(dataOut507) 
	 ,.R_out(R508) ,.data_out(dataOut508)  );
medianFilterCell  m509(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R508) ,.dataR_in(dataOut510) ,.dataL_in(dataOut508) 
	 ,.R_out(R509) ,.data_out(dataOut509)  );
medianFilterCell  m510(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R509) ,.dataR_in(dataOut511) ,.dataL_in(dataOut509) 
	 ,.R_out(R510) ,.data_out(dataOut510)  );
medianFilterCell  m511(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R510) ,.dataR_in(dataOut512) ,.dataL_in(dataOut510) 
	 ,.R_out(R511) ,.data_out(dataOut511)  );
medianFilterCell  m512(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R511) ,.dataR_in(dataOut513) ,.dataL_in(dataOut511) 
	 ,.R_out(R512) ,.data_out(dataOut512)  );
medianFilterCell  m513(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R512) ,.dataR_in(dataOut514) ,.dataL_in(dataOut512) 
	 ,.R_out(R513) ,.data_out(dataOut513)  );
medianFilterCell  m514(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R513) ,.dataR_in(dataOut515) ,.dataL_in(dataOut513) 
	 ,.R_out(R514) ,.data_out(dataOut514)  );
medianFilterCell  m515(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R514) ,.dataR_in(dataOut516) ,.dataL_in(dataOut514) 
	 ,.R_out(R515) ,.data_out(dataOut515)  );
medianFilterCell  m516(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R515) ,.dataR_in(dataOut517) ,.dataL_in(dataOut515) 
	 ,.R_out(R516) ,.data_out(dataOut516)  );
medianFilterCell  m517(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R516) ,.dataR_in(dataOut518) ,.dataL_in(dataOut516) 
	 ,.R_out(R517) ,.data_out(dataOut517)  );
medianFilterCell  m518(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R517) ,.dataR_in(dataOut519) ,.dataL_in(dataOut517) 
	 ,.R_out(R518) ,.data_out(dataOut518)  );
medianFilterCell  m519(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R518) ,.dataR_in(dataOut520) ,.dataL_in(dataOut518) 
	 ,.R_out(R519) ,.data_out(dataOut519)  );
medianFilterCell  m520(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R519) ,.dataR_in(dataOut521) ,.dataL_in(dataOut519) 
	 ,.R_out(R520) ,.data_out(dataOut520)  );
medianFilterCell  m521(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R520) ,.dataR_in(dataOut522) ,.dataL_in(dataOut520) 
	 ,.R_out(R521) ,.data_out(dataOut521)  );
medianFilterCell  m522(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R521) ,.dataR_in(dataOut523) ,.dataL_in(dataOut521) 
	 ,.R_out(R522) ,.data_out(dataOut522)  );
medianFilterCell  m523(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R522) ,.dataR_in(dataOut524) ,.dataL_in(dataOut522) 
	 ,.R_out(R523) ,.data_out(dataOut523)  );
medianFilterCell  m524(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R523) ,.dataR_in(dataOut525) ,.dataL_in(dataOut523) 
	 ,.R_out(R524) ,.data_out(dataOut524)  );
medianFilterCell  m525(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R524) ,.dataR_in(dataOut526) ,.dataL_in(dataOut524) 
	 ,.R_out(R525) ,.data_out(dataOut525)  );
medianFilterCell  m526(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R525) ,.dataR_in(dataOut527) ,.dataL_in(dataOut525) 
	 ,.R_out(R526) ,.data_out(dataOut526)  );
medianFilterCell  m527(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R526) ,.dataR_in(dataOut528) ,.dataL_in(dataOut526) 
	 ,.R_out(R527) ,.data_out(dataOut527)  );
medianFilterCell  m528(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R527) ,.dataR_in(dataOut529) ,.dataL_in(dataOut527) 
	 ,.R_out(R528) ,.data_out(dataOut528)  );
medianFilterCell  m529(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R528) ,.dataR_in(dataOut530) ,.dataL_in(dataOut528) 
	 ,.R_out(R529) ,.data_out(dataOut529)  );
medianFilterCell  m530(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R529) ,.dataR_in(dataOut531) ,.dataL_in(dataOut529) 
	 ,.R_out(R530) ,.data_out(dataOut530)  );
medianFilterCell  m531(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R530) ,.dataR_in(dataOut532) ,.dataL_in(dataOut530) 
	 ,.R_out(R531) ,.data_out(dataOut531)  );
medianFilterCell  m532(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R531) ,.dataR_in(dataOut533) ,.dataL_in(dataOut531) 
	 ,.R_out(R532) ,.data_out(dataOut532)  );
medianFilterCell  m533(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R532) ,.dataR_in(dataOut534) ,.dataL_in(dataOut532) 
	 ,.R_out(R533) ,.data_out(dataOut533)  );
medianFilterCell  m534(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R533) ,.dataR_in(dataOut535) ,.dataL_in(dataOut533) 
	 ,.R_out(R534) ,.data_out(dataOut534)  );
medianFilterCell  m535(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R534) ,.dataR_in(dataOut536) ,.dataL_in(dataOut534) 
	 ,.R_out(R535) ,.data_out(dataOut535)  );
medianFilterCell  m536(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R535) ,.dataR_in(dataOut537) ,.dataL_in(dataOut535) 
	 ,.R_out(R536) ,.data_out(dataOut536)  );
medianFilterCell  m537(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R536) ,.dataR_in(dataOut538) ,.dataL_in(dataOut536) 
	 ,.R_out(R537) ,.data_out(dataOut537)  );
medianFilterCell  m538(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R537) ,.dataR_in(dataOut539) ,.dataL_in(dataOut537) 
	 ,.R_out(R538) ,.data_out(dataOut538)  );
medianFilterCell  m539(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R538) ,.dataR_in(dataOut540) ,.dataL_in(dataOut538) 
	 ,.R_out(R539) ,.data_out(dataOut539)  );
medianFilterCell  m540(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R539) ,.dataR_in(dataOut541) ,.dataL_in(dataOut539) 
	 ,.R_out(R540) ,.data_out(dataOut540)  );
medianFilterCell  m541(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R540) ,.dataR_in(dataOut542) ,.dataL_in(dataOut540) 
	 ,.R_out(R541) ,.data_out(dataOut541)  );
medianFilterCell  m542(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R541) ,.dataR_in(dataOut543) ,.dataL_in(dataOut541) 
	 ,.R_out(R542) ,.data_out(dataOut542)  );
medianFilterCell  m543(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R542) ,.dataR_in(dataOut544) ,.dataL_in(dataOut542) 
	 ,.R_out(R543) ,.data_out(dataOut543)  );
medianFilterCell  m544(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R543) ,.dataR_in(dataOut545) ,.dataL_in(dataOut543) 
	 ,.R_out(R544) ,.data_out(dataOut544)  );
medianFilterCell  m545(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R544) ,.dataR_in(dataOut546) ,.dataL_in(dataOut544) 
	 ,.R_out(R545) ,.data_out(dataOut545)  );
medianFilterCell  m546(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R545) ,.dataR_in(dataOut547) ,.dataL_in(dataOut545) 
	 ,.R_out(R546) ,.data_out(dataOut546)  );
medianFilterCell  m547(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R546) ,.dataR_in(dataOut548) ,.dataL_in(dataOut546) 
	 ,.R_out(R547) ,.data_out(dataOut547)  );
medianFilterCell  m548(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R547) ,.dataR_in(dataOut549) ,.dataL_in(dataOut547) 
	 ,.R_out(R548) ,.data_out(dataOut548)  );
medianFilterCell  m549(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R548) ,.dataR_in(dataOut550) ,.dataL_in(dataOut548) 
	 ,.R_out(R549) ,.data_out(dataOut549)  );
medianFilterCell  m550(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R549) ,.dataR_in(dataOut551) ,.dataL_in(dataOut549) 
	 ,.R_out(R550) ,.data_out(dataOut550)  );
medianFilterCell  m551(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R550) ,.dataR_in(dataOut552) ,.dataL_in(dataOut550) 
	 ,.R_out(R551) ,.data_out(dataOut551)  );
medianFilterCell  m552(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R551) ,.dataR_in(dataOut553) ,.dataL_in(dataOut551) 
	 ,.R_out(R552) ,.data_out(dataOut552)  );
medianFilterCell  m553(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R552) ,.dataR_in(dataOut554) ,.dataL_in(dataOut552) 
	 ,.R_out(R553) ,.data_out(dataOut553)  );
medianFilterCell  m554(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R553) ,.dataR_in(dataOut555) ,.dataL_in(dataOut553) 
	 ,.R_out(R554) ,.data_out(dataOut554)  );
medianFilterCell  m555(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R554) ,.dataR_in(dataOut556) ,.dataL_in(dataOut554) 
	 ,.R_out(R555) ,.data_out(dataOut555)  );
medianFilterCell  m556(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R555) ,.dataR_in(dataOut557) ,.dataL_in(dataOut555) 
	 ,.R_out(R556) ,.data_out(dataOut556)  );
medianFilterCell  m557(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R556) ,.dataR_in(dataOut558) ,.dataL_in(dataOut556) 
	 ,.R_out(R557) ,.data_out(dataOut557)  );
medianFilterCell  m558(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R557) ,.dataR_in(dataOut559) ,.dataL_in(dataOut557) 
	 ,.R_out(R558) ,.data_out(dataOut558)  );
medianFilterCell  m559(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R558) ,.dataR_in(dataOut560) ,.dataL_in(dataOut558) 
	 ,.R_out(R559) ,.data_out(dataOut559)  );
medianFilterCell  m560(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R559) ,.dataR_in(dataOut561) ,.dataL_in(dataOut559) 
	 ,.R_out(R560) ,.data_out(dataOut560)  );
medianFilterCell  m561(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R560) ,.dataR_in(dataOut562) ,.dataL_in(dataOut560) 
	 ,.R_out(R561) ,.data_out(dataOut561)  );
medianFilterCell  m562(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R561) ,.dataR_in(dataOut563) ,.dataL_in(dataOut561) 
	 ,.R_out(R562) ,.data_out(dataOut562)  );
medianFilterCell  m563(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R562) ,.dataR_in(dataOut564) ,.dataL_in(dataOut562) 
	 ,.R_out(R563) ,.data_out(dataOut563)  );
medianFilterCell  m564(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R563) ,.dataR_in(dataOut565) ,.dataL_in(dataOut563) 
	 ,.R_out(R564) ,.data_out(dataOut564)  );
medianFilterCell  m565(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R564) ,.dataR_in(dataOut566) ,.dataL_in(dataOut564) 
	 ,.R_out(R565) ,.data_out(dataOut565)  );
medianFilterCell  m566(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R565) ,.dataR_in(dataOut567) ,.dataL_in(dataOut565) 
	 ,.R_out(R566) ,.data_out(dataOut566)  );
medianFilterCell  m567(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R566) ,.dataR_in(dataOut568) ,.dataL_in(dataOut566) 
	 ,.R_out(R567) ,.data_out(dataOut567)  );
medianFilterCell  m568(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R567) ,.dataR_in(dataOut569) ,.dataL_in(dataOut567) 
	 ,.R_out(R568) ,.data_out(dataOut568)  );
medianFilterCell  m569(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R568) ,.dataR_in(dataOut570) ,.dataL_in(dataOut568) 
	 ,.R_out(R569) ,.data_out(dataOut569)  );
medianFilterCell  m570(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R569) ,.dataR_in(dataOut571) ,.dataL_in(dataOut569) 
	 ,.R_out(R570) ,.data_out(dataOut570)  );
medianFilterCell  m571(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R570) ,.dataR_in(dataOut572) ,.dataL_in(dataOut570) 
	 ,.R_out(R571) ,.data_out(dataOut571)  );
medianFilterCell  m572(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R571) ,.dataR_in(dataOut573) ,.dataL_in(dataOut571) 
	 ,.R_out(R572) ,.data_out(dataOut572)  );
medianFilterCell  m573(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R572) ,.dataR_in(dataOut574) ,.dataL_in(dataOut572) 
	 ,.R_out(R573) ,.data_out(dataOut573)  );
medianFilterCell  m574(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R573) ,.dataR_in(dataOut575) ,.dataL_in(dataOut573) 
	 ,.R_out(R574) ,.data_out(dataOut574)  );
medianFilterCell  m575(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R574) ,.dataR_in(dataOut576) ,.dataL_in(dataOut574) 
	 ,.R_out(R575) ,.data_out(dataOut575)  );
medianFilterCell  m576(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R575) ,.dataR_in(dataOut577) ,.dataL_in(dataOut575) 
	 ,.R_out(R576) ,.data_out(dataOut576)  );
medianFilterCell  m577(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R576) ,.dataR_in(dataOut578) ,.dataL_in(dataOut576) 
	 ,.R_out(R577) ,.data_out(dataOut577)  );
medianFilterCell  m578(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R577) ,.dataR_in(dataOut579) ,.dataL_in(dataOut577) 
	 ,.R_out(R578) ,.data_out(dataOut578)  );
medianFilterCell  m579(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R578) ,.dataR_in(dataOut580) ,.dataL_in(dataOut578) 
	 ,.R_out(R579) ,.data_out(dataOut579)  );
medianFilterCell  m580(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R579) ,.dataR_in(dataOut581) ,.dataL_in(dataOut579) 
	 ,.R_out(R580) ,.data_out(dataOut580)  );
medianFilterCell  m581(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R580) ,.dataR_in(dataOut582) ,.dataL_in(dataOut580) 
	 ,.R_out(R581) ,.data_out(dataOut581)  );
medianFilterCell  m582(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R581) ,.dataR_in(dataOut583) ,.dataL_in(dataOut581) 
	 ,.R_out(R582) ,.data_out(dataOut582)  );
medianFilterCell  m583(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R582) ,.dataR_in(dataOut584) ,.dataL_in(dataOut582) 
	 ,.R_out(R583) ,.data_out(dataOut583)  );
medianFilterCell  m584(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R583) ,.dataR_in(dataOut585) ,.dataL_in(dataOut583) 
	 ,.R_out(R584) ,.data_out(dataOut584)  );
medianFilterCell  m585(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R584) ,.dataR_in(dataOut586) ,.dataL_in(dataOut584) 
	 ,.R_out(R585) ,.data_out(dataOut585)  );
medianFilterCell  m586(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R585) ,.dataR_in(dataOut587) ,.dataL_in(dataOut585) 
	 ,.R_out(R586) ,.data_out(dataOut586)  );
medianFilterCell  m587(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R586) ,.dataR_in(dataOut588) ,.dataL_in(dataOut586) 
	 ,.R_out(R587) ,.data_out(dataOut587)  );
medianFilterCell  m588(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R587) ,.dataR_in(dataOut589) ,.dataL_in(dataOut587) 
	 ,.R_out(R588) ,.data_out(dataOut588)  );
medianFilterCell  m589(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R588) ,.dataR_in(dataOut590) ,.dataL_in(dataOut588) 
	 ,.R_out(R589) ,.data_out(dataOut589)  );
medianFilterCell  m590(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R589) ,.dataR_in(dataOut591) ,.dataL_in(dataOut589) 
	 ,.R_out(R590) ,.data_out(dataOut590)  );
medianFilterCell  m591(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R590) ,.dataR_in(dataOut592) ,.dataL_in(dataOut590) 
	 ,.R_out(R591) ,.data_out(dataOut591)  );
medianFilterCell  m592(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R591) ,.dataR_in(dataOut593) ,.dataL_in(dataOut591) 
	 ,.R_out(R592) ,.data_out(dataOut592)  );
medianFilterCell  m593(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R592) ,.dataR_in(dataOut594) ,.dataL_in(dataOut592) 
	 ,.R_out(R593) ,.data_out(dataOut593)  );
medianFilterCell  m594(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R593) ,.dataR_in(dataOut595) ,.dataL_in(dataOut593) 
	 ,.R_out(R594) ,.data_out(dataOut594)  );
medianFilterCell  m595(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R594) ,.dataR_in(dataOut596) ,.dataL_in(dataOut594) 
	 ,.R_out(R595) ,.data_out(dataOut595)  );
medianFilterCell  m596(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R595) ,.dataR_in(dataOut597) ,.dataL_in(dataOut595) 
	 ,.R_out(R596) ,.data_out(dataOut596)  );
medianFilterCell  m597(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R596) ,.dataR_in(dataOut598) ,.dataL_in(dataOut596) 
	 ,.R_out(R597) ,.data_out(dataOut597)  );
medianFilterCell  m598(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R597) ,.dataR_in(dataOut599) ,.dataL_in(dataOut597) 
	 ,.R_out(R598) ,.data_out(dataOut598)  );
medianFilterCell  m599(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R598) ,.dataR_in(dataOut600) ,.dataL_in(dataOut598) 
	 ,.R_out(R599) ,.data_out(dataOut599)  );
medianFilterCell  m600(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R599) ,.dataR_in(dataOut601) ,.dataL_in(dataOut599) 
	 ,.R_out(R600) ,.data_out(dataOut600)  );
medianFilterCell  m601(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R600) ,.dataR_in(dataOut602) ,.dataL_in(dataOut600) 
	 ,.R_out(R601) ,.data_out(dataOut601)  );
medianFilterCell  m602(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R601) ,.dataR_in(dataOut603) ,.dataL_in(dataOut601) 
	 ,.R_out(R602) ,.data_out(dataOut602)  );
medianFilterCell  m603(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R602) ,.dataR_in(dataOut604) ,.dataL_in(dataOut602) 
	 ,.R_out(R603) ,.data_out(dataOut603)  );
medianFilterCell  m604(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R603) ,.dataR_in(dataOut605) ,.dataL_in(dataOut603) 
	 ,.R_out(R604) ,.data_out(dataOut604)  );
medianFilterCell  m605(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R604) ,.dataR_in(dataOut606) ,.dataL_in(dataOut604) 
	 ,.R_out(R605) ,.data_out(dataOut605)  );
medianFilterCell  m606(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R605) ,.dataR_in(dataOut607) ,.dataL_in(dataOut605) 
	 ,.R_out(R606) ,.data_out(dataOut606)  );
medianFilterCell  m607(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R606) ,.dataR_in(dataOut608) ,.dataL_in(dataOut606) 
	 ,.R_out(R607) ,.data_out(dataOut607)  );
medianFilterCell  m608(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R607) ,.dataR_in(dataOut609) ,.dataL_in(dataOut607) 
	 ,.R_out(R608) ,.data_out(dataOut608)  );
medianFilterCell  m609(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R608) ,.dataR_in(dataOut610) ,.dataL_in(dataOut608) 
	 ,.R_out(R609) ,.data_out(dataOut609)  );
medianFilterCell  m610(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R609) ,.dataR_in(dataOut611) ,.dataL_in(dataOut609) 
	 ,.R_out(R610) ,.data_out(dataOut610)  );
medianFilterCell  m611(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R610) ,.dataR_in(dataOut612) ,.dataL_in(dataOut610) 
	 ,.R_out(R611) ,.data_out(dataOut611)  );
medianFilterCell  m612(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R611) ,.dataR_in(dataOut613) ,.dataL_in(dataOut611) 
	 ,.R_out(R612) ,.data_out(dataOut612)  );
medianFilterCell  m613(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R612) ,.dataR_in(dataOut614) ,.dataL_in(dataOut612) 
	 ,.R_out(R613) ,.data_out(dataOut613)  );
medianFilterCell  m614(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R613) ,.dataR_in(dataOut615) ,.dataL_in(dataOut613) 
	 ,.R_out(R614) ,.data_out(dataOut614)  );
medianFilterCell  m615(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R614) ,.dataR_in(dataOut616) ,.dataL_in(dataOut614) 
	 ,.R_out(R615) ,.data_out(dataOut615)  );
medianFilterCell  m616(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R615) ,.dataR_in(dataOut617) ,.dataL_in(dataOut615) 
	 ,.R_out(R616) ,.data_out(dataOut616)  );
medianFilterCell  m617(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R616) ,.dataR_in(dataOut618) ,.dataL_in(dataOut616) 
	 ,.R_out(R617) ,.data_out(dataOut617)  );
medianFilterCell  m618(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R617) ,.dataR_in(dataOut619) ,.dataL_in(dataOut617) 
	 ,.R_out(R618) ,.data_out(dataOut618)  );
medianFilterCell  m619(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R618) ,.dataR_in(dataOut620) ,.dataL_in(dataOut618) 
	 ,.R_out(R619) ,.data_out(dataOut619)  );
medianFilterCell  m620(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R619) ,.dataR_in(dataOut621) ,.dataL_in(dataOut619) 
	 ,.R_out(R620) ,.data_out(dataOut620)  );
medianFilterCell  m621(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R620) ,.dataR_in(dataOut622) ,.dataL_in(dataOut620) 
	 ,.R_out(R621) ,.data_out(dataOut621)  );
medianFilterCell  m622(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R621) ,.dataR_in(dataOut623) ,.dataL_in(dataOut621) 
	 ,.R_out(R622) ,.data_out(dataOut622)  );
medianFilterCell  m623(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R622) ,.dataR_in(dataOut624) ,.dataL_in(dataOut622) 
	 ,.R_out(R623) ,.data_out(dataOut623)  );
medianFilterCell  m624(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R623) ,.dataR_in(dataOut625) ,.dataL_in(dataOut623) 
	 ,.R_out(R624) ,.data_out(dataOut624)  );
medianFilterCell  m625(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R624) ,.dataR_in(dataOut626) ,.dataL_in(dataOut624) 
	 ,.R_out(R625) ,.data_out(dataOut625)  );
medianFilterCell  m626(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R625) ,.dataR_in(dataOut627) ,.dataL_in(dataOut625) 
	 ,.R_out(R626) ,.data_out(dataOut626)  );
medianFilterCell  m627(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R626) ,.dataR_in(dataOut628) ,.dataL_in(dataOut626) 
	 ,.R_out(R627) ,.data_out(dataOut627)  );
medianFilterCell  m628(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R627) ,.dataR_in(dataOut629) ,.dataL_in(dataOut627) 
	 ,.R_out(R628) ,.data_out(dataOut628)  );
medianFilterCell  m629(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R628) ,.dataR_in(dataOut630) ,.dataL_in(dataOut628) 
	 ,.R_out(R629) ,.data_out(dataOut629)  );
medianFilterCell  m630(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R629) ,.dataR_in(dataOut631) ,.dataL_in(dataOut629) 
	 ,.R_out(R630) ,.data_out(dataOut630)  );
medianFilterCell  m631(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R630) ,.dataR_in(dataOut632) ,.dataL_in(dataOut630) 
	 ,.R_out(R631) ,.data_out(dataOut631)  );
medianFilterCell  m632(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R631) ,.dataR_in(dataOut633) ,.dataL_in(dataOut631) 
	 ,.R_out(R632) ,.data_out(dataOut632)  );
medianFilterCell  m633(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R632) ,.dataR_in(dataOut634) ,.dataL_in(dataOut632) 
	 ,.R_out(R633) ,.data_out(dataOut633)  );
medianFilterCell  m634(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R633) ,.dataR_in(dataOut635) ,.dataL_in(dataOut633) 
	 ,.R_out(R634) ,.data_out(dataOut634)  );
medianFilterCell  m635(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R634) ,.dataR_in(dataOut636) ,.dataL_in(dataOut634) 
	 ,.R_out(R635) ,.data_out(dataOut635)  );
medianFilterCell  m636(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R635) ,.dataR_in(dataOut637) ,.dataL_in(dataOut635) 
	 ,.R_out(R636) ,.data_out(dataOut636)  );
medianFilterCell  m637(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R636) ,.dataR_in(dataOut638) ,.dataL_in(dataOut636) 
	 ,.R_out(R637) ,.data_out(dataOut637)  );
medianFilterCell  m638(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R637) ,.dataR_in(dataOut639) ,.dataL_in(dataOut637) 
	 ,.R_out(R638) ,.data_out(dataOut638)  );
medianFilterCell  m639(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R638) ,.dataR_in(dataOut640) ,.dataL_in(dataOut638) 
	 ,.R_out(R639) ,.data_out(dataOut639)  );
medianFilterCell  m640(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R639) ,.dataR_in(dataOut641) ,.dataL_in(dataOut639) 
	 ,.R_out(R640) ,.data_out(dataOut640)  );
medianFilterCell  m641(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R640) ,.dataR_in(dataOut642) ,.dataL_in(dataOut640) 
	 ,.R_out(R641) ,.data_out(dataOut641)  );
medianFilterCell  m642(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R641) ,.dataR_in(dataOut643) ,.dataL_in(dataOut641) 
	 ,.R_out(R642) ,.data_out(dataOut642)  );
medianFilterCell  m643(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R642) ,.dataR_in(dataOut644) ,.dataL_in(dataOut642) 
	 ,.R_out(R643) ,.data_out(dataOut643)  );
medianFilterCell  m644(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R643) ,.dataR_in(dataOut645) ,.dataL_in(dataOut643) 
	 ,.R_out(R644) ,.data_out(dataOut644)  );
medianFilterCell  m645(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R644) ,.dataR_in(dataOut646) ,.dataL_in(dataOut644) 
	 ,.R_out(R645) ,.data_out(dataOut645)  );
medianFilterCell  m646(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R645) ,.dataR_in(dataOut647) ,.dataL_in(dataOut645) 
	 ,.R_out(R646) ,.data_out(dataOut646)  );
medianFilterCell  m647(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R646) ,.dataR_in(dataOut648) ,.dataL_in(dataOut646) 
	 ,.R_out(R647) ,.data_out(dataOut647)  );
medianFilterCell  m648(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R647) ,.dataR_in(dataOut649) ,.dataL_in(dataOut647) 
	 ,.R_out(R648) ,.data_out(dataOut648)  );
medianFilterCell  m649(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R648) ,.dataR_in(dataOut650) ,.dataL_in(dataOut648) 
	 ,.R_out(R649) ,.data_out(dataOut649)  );
medianFilterCell  m650(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R649) ,.dataR_in(dataOut651) ,.dataL_in(dataOut649) 
	 ,.R_out(R650) ,.data_out(dataOut650)  );
medianFilterCell  m651(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R650) ,.dataR_in(dataOut652) ,.dataL_in(dataOut650) 
	 ,.R_out(R651) ,.data_out(dataOut651)  );
medianFilterCell  m652(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R651) ,.dataR_in(dataOut653) ,.dataL_in(dataOut651) 
	 ,.R_out(R652) ,.data_out(dataOut652)  );
medianFilterCell  m653(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R652) ,.dataR_in(dataOut654) ,.dataL_in(dataOut652) 
	 ,.R_out(R653) ,.data_out(dataOut653)  );
medianFilterCell  m654(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R653) ,.dataR_in(dataOut655) ,.dataL_in(dataOut653) 
	 ,.R_out(R654) ,.data_out(dataOut654)  );
medianFilterCell  m655(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R654) ,.dataR_in(dataOut656) ,.dataL_in(dataOut654) 
	 ,.R_out(R655) ,.data_out(dataOut655)  );
medianFilterCell  m656(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R655) ,.dataR_in(dataOut657) ,.dataL_in(dataOut655) 
	 ,.R_out(R656) ,.data_out(dataOut656)  );
medianFilterCell  m657(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R656) ,.dataR_in(dataOut658) ,.dataL_in(dataOut656) 
	 ,.R_out(R657) ,.data_out(dataOut657)  );
medianFilterCell  m658(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R657) ,.dataR_in(dataOut659) ,.dataL_in(dataOut657) 
	 ,.R_out(R658) ,.data_out(dataOut658)  );
medianFilterCell  m659(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R658) ,.dataR_in(dataOut660) ,.dataL_in(dataOut658) 
	 ,.R_out(R659) ,.data_out(dataOut659)  );
medianFilterCell  m660(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R659) ,.dataR_in(dataOut661) ,.dataL_in(dataOut659) 
	 ,.R_out(R660) ,.data_out(dataOut660)  );
medianFilterCell  m661(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R660) ,.dataR_in(dataOut662) ,.dataL_in(dataOut660) 
	 ,.R_out(R661) ,.data_out(dataOut661)  );
medianFilterCell  m662(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R661) ,.dataR_in(dataOut663) ,.dataL_in(dataOut661) 
	 ,.R_out(R662) ,.data_out(dataOut662)  );
medianFilterCell  m663(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R662) ,.dataR_in(dataOut664) ,.dataL_in(dataOut662) 
	 ,.R_out(R663) ,.data_out(dataOut663)  );
medianFilterCell  m664(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R663) ,.dataR_in(dataOut665) ,.dataL_in(dataOut663) 
	 ,.R_out(R664) ,.data_out(dataOut664)  );
medianFilterCell  m665(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R664) ,.dataR_in(dataOut666) ,.dataL_in(dataOut664) 
	 ,.R_out(R665) ,.data_out(dataOut665)  );
medianFilterCell  m666(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R665) ,.dataR_in(dataOut667) ,.dataL_in(dataOut665) 
	 ,.R_out(R666) ,.data_out(dataOut666)  );
medianFilterCell  m667(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R666) ,.dataR_in(dataOut668) ,.dataL_in(dataOut666) 
	 ,.R_out(R667) ,.data_out(dataOut667)  );
medianFilterCell  m668(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R667) ,.dataR_in(dataOut669) ,.dataL_in(dataOut667) 
	 ,.R_out(R668) ,.data_out(dataOut668)  );
medianFilterCell  m669(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R668) ,.dataR_in(dataOut670) ,.dataL_in(dataOut668) 
	 ,.R_out(R669) ,.data_out(dataOut669)  );
medianFilterCell  m670(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R669) ,.dataR_in(dataOut671) ,.dataL_in(dataOut669) 
	 ,.R_out(R670) ,.data_out(dataOut670)  );
medianFilterCell  m671(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R670) ,.dataR_in(dataOut672) ,.dataL_in(dataOut670) 
	 ,.R_out(R671) ,.data_out(dataOut671)  );
medianFilterCell  m672(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R671) ,.dataR_in(dataOut673) ,.dataL_in(dataOut671) 
	 ,.R_out(R672) ,.data_out(dataOut672)  );
medianFilterCell  m673(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R672) ,.dataR_in(dataOut674) ,.dataL_in(dataOut672) 
	 ,.R_out(R673) ,.data_out(dataOut673)  );
medianFilterCell  m674(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R673) ,.dataR_in(dataOut675) ,.dataL_in(dataOut673) 
	 ,.R_out(R674) ,.data_out(dataOut674)  );
medianFilterCell  m675(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R674) ,.dataR_in(dataOut676) ,.dataL_in(dataOut674) 
	 ,.R_out(R675) ,.data_out(dataOut675)  );
medianFilterCell  m676(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R675) ,.dataR_in(dataOut677) ,.dataL_in(dataOut675) 
	 ,.R_out(R676) ,.data_out(dataOut676)  );
medianFilterCell  m677(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R676) ,.dataR_in(dataOut678) ,.dataL_in(dataOut676) 
	 ,.R_out(R677) ,.data_out(dataOut677)  );
medianFilterCell  m678(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R677) ,.dataR_in(dataOut679) ,.dataL_in(dataOut677) 
	 ,.R_out(R678) ,.data_out(dataOut678)  );
medianFilterCell  m679(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R678) ,.dataR_in(dataOut680) ,.dataL_in(dataOut678) 
	 ,.R_out(R679) ,.data_out(dataOut679)  );
medianFilterCell  m680(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R679) ,.dataR_in(dataOut681) ,.dataL_in(dataOut679) 
	 ,.R_out(R680) ,.data_out(dataOut680)  );
medianFilterCell  m681(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R680) ,.dataR_in(dataOut682) ,.dataL_in(dataOut680) 
	 ,.R_out(R681) ,.data_out(dataOut681)  );
medianFilterCell  m682(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R681) ,.dataR_in(dataOut683) ,.dataL_in(dataOut681) 
	 ,.R_out(R682) ,.data_out(dataOut682)  );
medianFilterCell  m683(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R682) ,.dataR_in(dataOut684) ,.dataL_in(dataOut682) 
	 ,.R_out(R683) ,.data_out(dataOut683)  );
medianFilterCell  m684(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R683) ,.dataR_in(dataOut685) ,.dataL_in(dataOut683) 
	 ,.R_out(R684) ,.data_out(dataOut684)  );
medianFilterCell  m685(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R684) ,.dataR_in(dataOut686) ,.dataL_in(dataOut684) 
	 ,.R_out(R685) ,.data_out(dataOut685)  );
medianFilterCell  m686(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R685) ,.dataR_in(dataOut687) ,.dataL_in(dataOut685) 
	 ,.R_out(R686) ,.data_out(dataOut686)  );
medianFilterCell  m687(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R686) ,.dataR_in(dataOut688) ,.dataL_in(dataOut686) 
	 ,.R_out(R687) ,.data_out(dataOut687)  );
medianFilterCell  m688(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R687) ,.dataR_in(dataOut689) ,.dataL_in(dataOut687) 
	 ,.R_out(R688) ,.data_out(dataOut688)  );
medianFilterCell  m689(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R688) ,.dataR_in(dataOut690) ,.dataL_in(dataOut688) 
	 ,.R_out(R689) ,.data_out(dataOut689)  );
medianFilterCell  m690(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R689) ,.dataR_in(dataOut691) ,.dataL_in(dataOut689) 
	 ,.R_out(R690) ,.data_out(dataOut690)  );
medianFilterCell  m691(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R690) ,.dataR_in(dataOut692) ,.dataL_in(dataOut690) 
	 ,.R_out(R691) ,.data_out(dataOut691)  );
medianFilterCell  m692(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R691) ,.dataR_in(dataOut693) ,.dataL_in(dataOut691) 
	 ,.R_out(R692) ,.data_out(dataOut692)  );
medianFilterCell  m693(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R692) ,.dataR_in(dataOut694) ,.dataL_in(dataOut692) 
	 ,.R_out(R693) ,.data_out(dataOut693)  );
medianFilterCell  m694(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R693) ,.dataR_in(dataOut695) ,.dataL_in(dataOut693) 
	 ,.R_out(R694) ,.data_out(dataOut694)  );
medianFilterCell  m695(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R694) ,.dataR_in(dataOut696) ,.dataL_in(dataOut694) 
	 ,.R_out(R695) ,.data_out(dataOut695)  );
medianFilterCell  m696(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R695) ,.dataR_in(dataOut697) ,.dataL_in(dataOut695) 
	 ,.R_out(R696) ,.data_out(dataOut696)  );
medianFilterCell  m697(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R696) ,.dataR_in(dataOut698) ,.dataL_in(dataOut696) 
	 ,.R_out(R697) ,.data_out(dataOut697)  );
medianFilterCell  m698(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R697) ,.dataR_in(dataOut699) ,.dataL_in(dataOut697) 
	 ,.R_out(R698) ,.data_out(dataOut698)  );
medianFilterCell  m699(.X(X) ,.oldData(oldData)  ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R698) ,.dataR_in(dataOut700) ,.dataL_in(dataOut698) 
	 ,.R_out(R699) ,.data_out(dataOut699)  );
medianFilterCell  m700(.X(X) ,.oldData(oldData) ,.flag(flag),.reset(reset) ,.clk(clk) ,.R_in(R699),.dataR_in(0) ,.dataL_in(dataOut699) 
	 ,.R_out(R700)  ,.data_out(dataOut700));


endmodule